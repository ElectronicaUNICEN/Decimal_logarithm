-- el resultado <ln> est� normalizado en 0.yyyyyyy (para precisi�n 7)
-- en 0.yyyyyyyyyyyyyyyy (para precisi�n 16)
-- en 0.yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy (para precisi�n 34)

-- cuando step es igual a 1, algunas celdas LUTS(1) no sopn usadas, ya que se opero de modo que 0.7<=x(1)<1.4

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.my_package.all;

Library UNISIM;
use UNISIM.vcomponents.all;

entity Lut_log is
	generic (P: integer:=7);
    port ( step : in  STD_LOGIC_VECTOR (log2sup(P)-1 downto 0); 
           d : in  STD_LOGIC_VECTOR (3 downto 0);-- corresponde a xi
			  step_eq_0: in std_logic; -- indica si step es igual a 0
			  x_greater_1: in std_logic; -- infdica si x es mayor a uno
           log : out  STD_LOGIC_VECTOR (4*P downto 0)); -- en SVA, por eso un bit m�s
end Lut_log;


architecture Behavioral of Lut_log is


-- == Comienzo declaraci�n
-- =============== Memoria LUT correspondiente a los ln c(i), usado solo en step=0 


type mlut_Log_0 is array (0 to 9) of std_logic_vector (4*P-1 downto 0);
---- los resultados est�n normalizados en 0.yyyyyyy (para precisi�n 7),
---- en 0.yyyyyyyyyyyyyyyy (para precisi�n 16)
---- en 0.yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy (para precisi�n 34)
--
signal lut_Log: mlut_Log_0 := ( 
		x"0000000", -- LUT(0), No usada
		x"8450980", -- LUT(1), ln 7 = 0.84509804001425683071221625859264
		x"6020599", -- LUT(2), ln 4 = 0.60205999132796239042747778944899
		x"4771212", -- LUT(3), ln 3 = 0.47712125471966243729502790325512
		x"3010299", -- LUT(4), ln 2 = 0.30102999566398119521373889472449
		x"3010299", -- LUT(5), ln 2 = 0.30102999566398119521373889472449
		x"3010299", -- LUT(6), ln 2 = 0.30102999566398119521373889472449
		x"0000000", -- LUT(7), ln 1 = 0.000000
		x"0000000", -- LUT(8), ln 1 = 0.000000
		x"0000000"); -- LUT(9), ln 1 = 0.000000



--signal lut_Log: mlut_Log_0 := ( 
--		x"0000000000000000", -- LUT(0), No usada
--		x"8450980400142568", -- LUT(1), ln 7 = 0.84509804001425683071221625859264
--		x"6020599913279623", -- LUT(2), ln 4 = 0.60205999132796239042747778944899
--		x"4771212547196624", -- LUT(3), ln 3 = 0.47712125471966243729502790325512
--		x"3010299956639811", -- LUT(4), ln 2 = 0.30102999566398119521373889472449
--		x"3010299956639811", -- LUT(5), ln 2 = 0.30102999566398119521373889472449
--		x"3010299956639811", -- LUT(6), ln 2 = 0.30102999566398119521373889472449
--		x"0000000000000000", -- LUT(7), ln 1 = 0.000000
--		x"0000000000000000", -- LUT(8), ln 1 = 0.000000
--		x"0000000000000000"); -- LUT(9), ln 1 = 0.000000

----
--signal lut_Log: mlut_Log_0 := ( 
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"8450980400142568307122162585926400", -- LUT(1), ln 7 = 0.84509804001425683071221625859264
--		x"6020599913279623904274777894489900", -- LUT(2), ln 4 = 0.60205999132796239042747778944899
--		x"4771212547196624372950279032551200", -- LUT(3), ln 3 = 0.47712125471966243729502790325512
--		x"3010299956639811952137388947244900", -- LUT(4), ln 2 = 0.30102999566398119521373889472449
--		x"3010299956639811952137388947244900", -- LUT(5), ln 2 = 0.30102999566398119521373889472449
--		x"3010299956639811952137388947244900", -- LUT(6), ln 2 = 0.30102999566398119521373889472449
--		x"0000000000000000000000000000000000", -- LUT(7), ln 1 = 0.000000
--		x"0000000000000000000000000000000000", -- LUT(8), ln 1 = 0.000000
--		x"0000000000000000000000000000000000"); -- LUT(9), ln 1 = 0.000000

	
-- ====== Comienzo declaraci�n
-- declaracion de meomria de ln para la parte de x>1

type mlut_LogShP is array (0 to P-1) of std_logic_vector (4*P-1 downto 0);
-- los resultados est�n normalizados en 0.yyyyyyy (para precisi�n 7),
-- en 0.yyyyyyyyyyyyyyyy (para precisi�n 16)
-- en 0.yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy (para precisi�n 34)

signal lut_Log10ShP1: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"0457574", -- LUT(1) = log10 (0.9) = -0.045757491
		x"0043648", -- LUT(2) = log10 (0.99) = -0.0043648054
		x"0004345", -- LUT(3) = log10 (0.999) = -0.00043451177
		x"0000434", -- LUT(4) = log10 (0.9999) = -0.000043431620
		x"0000043", -- LUT(5) = log10 (0.99999) = -0.0000043429665
		x"0000004"); -- LUT(6) = log10 (0.999999) = -4.3429470E-7

signal lut_Log10ShP2: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"0969100", -- LUT(1) = log10 (0.8) = -0.096910013
		x"0087739", -- LUT(2) = log10 (0.98) = -0.0087739243
		x"0008694", -- LUT(3) = log10 (0.998) = -0.00086945871
		x"0000868", -- LUT(4) = log10 (0.9998) = -0.000086867583
		x"0000086", -- LUT(5) = log10 (0.99998) = -0.0000086859765
		x"0000008"); -- LUT(6) = log10 (0.999998) = -8.6858983E-7

signal lut_Log10ShP3: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"1549019", -- LUT(1) = log10 (0.7) = -0.15490196
		x"0132282", -- LUT(2) = log10 (0.97) = -0.013228266
		x"0013048", -- LUT(3) = log10 (0.997) = -0.0013048417
		x"0001303", -- LUT(4) = log10 (0.9997) = -0.00013030789
		x"0000130", -- LUT(5) = log10 (0.99997) = -0.000013029030
		x"0000013"); -- LUT(6) = log10 (0.999997) = -0.0000013028854

signal lut_Log10ShP4: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"2218487", -- LUT(1) = log10 (0.6) = -0.22184875
		x"0177287", -- LUT(2) = log10 (0.96) = -0.017728767
		x"0017406", -- LUT(3) = log10 (0.996) = -0.0017406616
		x"0001737", -- LUT(4) = log10 (0.9996) = -0.00017375255
		x"0000173", -- LUT(5) = log10 (0.99996) = -0.000017372127
		x"0000017"); -- LUT(6) = log10 (0.999996) = -0.0000017371814

signal lut_Log10ShP5: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"3010300", -- LUT(1) = log10 (0.5) = -0.30103000
		x"0222763", -- LUT(2) = log10 (0.95) = -0.022276395
		x"0021769", -- LUT(3) = log10 (0.995) = -0.0021769193
		x"0002172", -- LUT(4) = log10 (0.9995) = -0.00021720155
		x"0000217", -- LUT(5) = log10 (0.99995) = -0.000021715267
		x"0000021"); -- LUT(6) = log10 (0.999995) = -0.0000021714778

signal lut_Log10ShP6: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"3979400", -- LUT(1) = log10 (0.4) = -0.39794001
		x"0268721", -- LUT(2) = log10 (0.94) = -0.026872146
		x"0026136", -- LUT(3) = log10 (0.994) = -0.0026136156
		x"0002606", -- LUT(4) = log10 (0.9994) = -0.00026065489
		x"0000260", -- LUT(5) = log10 (0.99994) = -0.000026058451
		x"0000026"); -- LUT(6) = log10 (0.999994) = -0.0000026057747

signal lut_Log10ShP7: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"5228787", -- LUT(1) = log10 (0.3) = -0.52287875
		x"0315170", -- LUT(2) = log10 (0.93) = -0.031517051
		x"0030507", -- LUT(3) = log10 (0.993) = -0.0030507515
		x"0003041", -- LUT(4) = log10 (0.9993) = -0.00030411259
		x"0000304", -- LUT(5) = log10 (0.99993) = -0.000030401678
		x"0000030"); -- LUT(6) = log10 (0.999993) = -0.0000030400720

signal lut_Log10ShP8: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"6989700", -- LUT(1) = log10 (0.2) = -0.69897000
		x"0362121", -- LUT(2) = log10 (0.92) = -0.036212173
		x"0034883", -- LUT(3) = log10 (0.992) = -0.0034883278
		x"0003475", -- LUT(4) = log10 (0.9992) = -0.00034757463
		x"0000347", -- LUT(5) = log10 (0.99992) = -0.000034744948
		x"0000034"); -- LUT(6) = log10 (0.999992) = -0.0000034743698

signal lut_Log10ShP9: mlut_LogShP := (
		x"0000000", -- LUT(0), No usada
		x"0000000", -- LUT(1) = log10 (0.1) = -1
		x"0409586", -- LUT(2) = log10 (0.91) = -0.040958608
		x"0039263", -- LUT(3) = log10 (0.991) = -0.0039263455
		x"0003910", -- LUT(4) = log10 (0.9991) = -0.00039104103
		x"0000390", -- LUT(5) = log10 (0.99991) = -0.000039088262
		x"0000039"); -- LUT(6) = log10 (0.999991) = -0.0000039086679
--
--signal lut_Log10ShP1: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"0457574905606751", -- LUT(1) = log10 (0.9) = -0.045757490560675125
--		x"0043648054024500", -- LUT(2) = log10 (0.99) = -0.0043648054024500847
--		x"0004345117740176", -- LUT(3) = log10 (0.999) = -0.00043451177401769131
--		x"0000434316198075", -- LUT(4) = log10 (0.9999) = -0.000043431619807510385
--		x"0000043429665339", -- LUT(5) = log10 (0.99999) = -0.0000043429665339013794
--		x"0000004342946990", -- LUT(6) = log10 (0.999999) = -4.3429469905063754E-7
--		x"0000000434294503", -- LUT(7) = log10 (0.9999999) = -4.3429450361797737E-8
--		x"0000000043429448", -- LUT(8) = log10 (0.99999999) = -4.3429448407472425E-9
--		x"0000000004342944", -- LUT(9) = log10 (0.999999999) = -4.3429448212039907E-10
--		x"0000000000434294", -- LUT(10) = log10 (0.9999999999) = -4.3429448192496655E-11
--		x"0000000000043429", -- LUT(11) = log10 (0.99999999999) = -4.3429448190542330E-12
--		x"0000000000004342", -- LUT(12) = log10 (0.999999999999) = -4.3429448190346897E-13
--		x"0000000000000434", -- LUT(13) = log10 (0.9999999999999) = -4.3429448190327354E-14
--		x"0000000000000043", -- LUT(14) = log10 (0.99999999999999) = -4.3429448190325400E-15
--		x"0000000000000004"); -- LUT(15) = log10 (0.999999999999999) = -4.3429448190325204E-16
--
--
--
--signal lut_Log10ShP2: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"0969100130080564", -- LUT(1) = log10 (0.8) = -0.096910013008056414
--		x"0087739243075051", -- LUT(2) = log10 (0.98) = -0.0087739243075051434
--		x"0008694587126288", -- LUT(3) = log10 (0.998) = -0.00086945871262889062
--		x"0000868675834285", -- LUT(4) = log10 (0.9998) = -0.000086867583428580795
--		x"0000086859764981", -- LUT(5) = log10 (0.99998) = -0.0000086859764981195532
--		x"0000008685898323", -- LUT(6) = log10 (0.999998) = -8.6858983239662558E-7
--		x"0000000868589050", -- LUT(7) = log10 (0.9999998) = -8.6858905066541162E-8
--		x"0000000086858897", -- LUT(8) = log10 (0.99999998) = -8.6858897249239341E-9
--		x"0000000008685889", -- LUT(9) = log10 (0.999999998) = -8.6858896467509262E-10
--		x"0000000000868588", -- LUT(10) = log10 (0.9999999998) = -8.6858896389336255E-11
--		x"0000000000086858", -- LUT(11) = log10 (0.99999999998) = -8.6858896381518954E-12
--		x"0000000000008685", -- LUT(12) = log10 (0.999999999998) = -8.6858896380737224E-13
--		x"0000000000000868", -- LUT(13) = log10 (0.9999999999998) = -8.6858896380659051E-14
--		x"0000000000000086", -- LUT(14) = log10 (0.99999999999998) = -8.6858896380651234E-15
--		x"0000000000000008"); -- LUT(15) = log10 (0.999999999999998) = -8.6858896380650452E-16
--
--signal lut_Log10ShP3: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"1549019599857431", -- LUT(1) = log10 (0.7) = -0.15490195998574317
--		x"0132282657337551", -- LUT(2) = log10 (0.97) = -0.013228265733755148
--		x"0013048416883442", -- LUT(3) = log10 (0.997) = -0.0013048416883442801
--		x"0001303078917321", -- LUT(4) = log10 (0.9997) = -0.00013030789173219119
--		x"0000130290298935", -- LUT(5) = log10 (0.99997) = -0.000013029029893523150
--		x"0000013028854000", -- LUT(6) = log10 (0.999997) = -0.0000013028854000388327
--		x"0000001302883641", -- LUT(7) = log10 (0.9999997) = -1.3028836411423114E-7
--		x"0000000130288346", -- LUT(8) = log10 (0.99999997) = -1.3028834652530076E-8
--		x"0000000013028834", -- LUT(9) = log10 (0.999999997) = -1.3028834476640807E-9
--		x"0000000001302883", -- LUT(10) = log10 (0.9999999997) = -1.3028834459051880E-10
--		x"0000000000130288", -- LUT(11) = log10 (0.99999999997) = -1.3028834457292987E-11
--		x"0000000000013028", -- LUT(12) = log10 (0.999999999997) = -1.3028834457117098E-12
--		x"0000000000001302", -- LUT(13) = log10 (0.9999999999997) = -1.3028834457099509E-13
--		x"0000000000000130", -- LUT(14) = log10 (0.99999999999997) = -1.3028834457097750E-14
--		x"0000000000000013"); -- LUT(15) = log10 (0.999999999999997) = -1.3028834457097574E-15
--
--signal lut_Log10ShP4: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"2218487496163563", -- LUT(1) = log10 (0.6) = -0.22184874961635637
--		x"0177287669604315", -- LUT(2) = log10 (0.96) = -0.017728766960431587
--		x"0017406615763012", -- LUT(3) = log10 (0.996) = -0.0017406615763012684
--		x"0001737525455875", -- LUT(4) = log10 (0.9996) = -0.00017375254558758231
--		x"0000173721267209", -- LUT(5) = log10 (0.99996) = -0.000017372126720980823
--		x"0000017371814019", -- LUT(6) = log10 (0.999996) = -0.0000017371814019781275
--		x"0000001737178275", -- LUT(7) = log10 (0.9999996) = -1.7371782750486855E-7
--		x"0000000173717796", -- LUT(8) = log10 (0.99999996) = -1.7371779623565668E-8
--		x"0000000017371779", -- LUT(9) = log10 (0.999999996) = -1.7371779310873632E-9
--		x"0000000001737177", -- LUT(10) = log10 (0.9999999996) = -1.7371779279604429E-10
--		x"0000000000173717", -- LUT(11) = log10 (0.99999999996) = -1.7371779276477509E-11
--		x"0000000000017371", -- LUT(12) = log10 (0.999999999996) = -1.7371779276164817E-12
--		x"0000000000001737", -- LUT(13) = log10 (0.9999999999996) = -1.7371779276133547E-13
--		x"0000000000000173", -- LUT(14) = log10 (0.99999999999996) = -1.7371779276130421E-14
--		x"0000000000000017"); -- LUT(15) = log10 (0.999999999999996) = -1.7371779276130108E-15
--
--signal lut_Log10ShP5: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"3010299956639812", -- LUT(1) = log10 (0.5) = -0.30102999566398120
--		x"0222763947111522", -- LUT(2) = log10 (0.95) = -0.022276394711152234
--		x"0021769192542745", -- LUT(3) = log10 (0.995) = -0.0021769192542745451
--		x"0002172015458642", -- LUT(4) = log10 (0.9995) = -0.00021720154586425580
--		x"0000217152669813", -- LUT(5) = log10 (0.99995) = -0.000021715266981361252
--		x"0000021714778382", -- LUT(6) = log10 (0.999995) = -0.0000021714778382153786
--		x"0000002171472952", -- LUT(7) = log10 (0.9999995) = -2.1714729523845425E-7
--		x"0000000217147246", -- LUT(8) = log10 (0.99999995) = -2.1714724638030712E-8
--		x"0000000021714724", -- LUT(9) = log10 (0.999999995) = -2.1714724149449402E-9
--		x"0000000002171472", -- LUT(10) = log10 (0.9999999995) = -2.1714724100591272E-10
--		x"0000000000217147", -- LUT(11) = log10 (0.99999999995) = -2.1714724095705459E-11
--		x"0000000000021714", -- LUT(12) = log10 (0.999999999995) = -2.1714724095216878E-12
--		x"0000000000002171", -- LUT(13) = log10 (0.9999999999995) = -2.1714724095168020E-13
--		x"0000000000000217", -- LUT(14) = log10 (0.99999999999995) = -2.1714724095163134E-14
--		x"0000000000000021"); -- LUT(15) = log10 (0.999999999999995) = -2.1714724095162646E-15
--
--signal lut_Log10ShP6: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"3979400086720376", -- LUT(1) = log10 (0.4) = -0.39794000867203761
--		x"0268721464003013", -- LUT(2) = log10 (0.94) = -0.026872146400301340
--		x"0026136156026866", -- LUT(3) = log10 (0.994) = -0.0026136156026866880
--		x"0002606548934319", -- LUT(4) = log10 (0.9994) = -0.00026065489343197428
--		x"0000260584506755", -- LUT(5) = log10 (0.99994) = -0.000026058450675533145
--		x"0000026057747087", -- LUT(6) = log10 (0.999994) = -0.0000026057747087514546
--		x"0000002605767673", -- LUT(7) = log10 (0.9999994) = -2.6057676731498911E-7
--		x"0000000260576696", -- LUT(8) = log10 (0.99999994) = -2.6057669695925208E-8
--		x"0000000026057668", -- LUT(9) = log10 (0.999999994) = -2.6057668992368117E-9
--		x"0000000002605766", -- LUT(10) = log10 (0.9999999994) = -2.6057668922012410E-10
--		x"0000000000260576", -- LUT(11) = log10 (0.99999999994) = -2.6057668914976840E-11
--		x"0000000000026057", -- LUT(12) = log10 (0.999999999994) = -2.6057668914273283E-12
--		x"0000000000002605", -- LUT(13) = log10 (0.9999999999994) = -2.6057668914202927E-13
--		x"0000000000000260", -- LUT(14) = log10 (0.99999999999994) = -2.6057668914195891E-14
--		x"0000000000000026"); -- LUT(15) = log10 (0.999999999999994) = -2.6057668914195188E-15
--
--signal lut_Log10ShP7: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"5228787452803375", -- LUT(1) = log10 (0.3) = -0.52287874528033756
--		x"0315170514460648", -- LUT(2) = log10 (0.93) = -0.031517051446064883
--		x"0030507515046188", -- LUT(3) = log10 (0.993) = -0.0030507515046188241
--		x"0003041125891607", -- LUT(4) = log10 (0.9993) = -0.00030411258916076147
--		x"0000304016778043", -- LUT(5) = log10 (0.99993) = -0.000030401677804365234
--		x"0000030400720135", -- LUT(6) = log10 (0.999993) = -0.0000030400720135872240
--		x"0000003040062437", -- LUT(7) = log10 (0.9999993) = -3.0400624373447400E-7
--		x"0000000304006147", -- LUT(8) = log10 (0.99999993) = -3.0400614797249158E-8
--		x"0000000030400613", -- LUT(9) = log10 (0.999999993) = -3.0400613839629776E-9
--		x"0000000003040061", -- LUT(10) = log10 (0.9999999993) = -3.0400613743867843E-10
--		x"0000000000304006", -- LUT(11) = log10 (0.99999999993) = -3.0400613734291649E-11
--		x"0000000000030400", -- LUT(12) = log10 (0.999999999993) = -3.0400613733334030E-12
--		x"0000000000003040", -- LUT(13) = log10 (0.9999999999993) = -3.0400613733238268E-13
--		x"0000000000000304", -- LUT(14) = log10 (0.99999999999993) = -3.0400613733228692E-14
--		x"0000000000000030"); -- LUT(15) = log10 (0.999999999999993) = -3.0400613733227734E-15
--
--signal lut_Log10ShP8: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"6989700043360188", -- LUT(1) = log10 (0.2) = -0.69897000433601880
--		x"0362121726544447", -- LUT(2) = log10 (0.92) = -0.036212172654444731
--		x"0034883278458213", -- LUT(3) = log10 (0.992) = -0.0034883278458213443
--		x"0003475746339209", -- LUT(4) = log10 (0.9992) = -0.00034757463392090232
--		x"0000347449483687", -- LUT(5) = log10 (0.99992) = -0.000034744948368726276
--		x"0000034743697527", -- LUT(6) = log10 (0.999992) = -0.0000034743697527235556
--		x"0000003474357244", -- LUT(7) = log10 (0.9999992) = -3.4743572449690979E-7
--		x"0000000347435599", -- LUT(8) = log10 (0.99999992) = -3.4743559942002562E-8
--		x"0000000034743558", -- LUT(9) = log10 (0.999999992) = -3.4743558691234381E-9
--		x"0000000003474355", -- LUT(10) = log10 (0.9999999992) = -3.4743558566157570E-10
--		x"0000000000347435", -- LUT(11) = log10 (0.99999999992) = -3.4743558553649889E-11
--		x"0000000000034743", -- LUT(12) = log10 (0.999999999992) = -3.4743558552399120E-12
--		x"0000000000003474", -- LUT(13) = log10 (0.9999999999992) = -3.4743558552274044E-13
--		x"0000000000000347", -- LUT(14) = log10 (0.99999999999992) = -3.4743558552261536E-14
--		x"0000000000000034"); -- LUT(15) = log10 (0.999999999999992) = -3.4743558552260285E-15
--
--signal lut_Log10ShP9: mlut_LogShP := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"0000000000000000", -- LUT(1) = log10 (0.1) = -1
--		x"0409586076789064", -- LUT(2) = log10 (0.91) = -0.040958607678906400
--		x"0039263455147246", -- LUT(3) = log10 (0.991) = -0.0039263455147246716
--		x"0003910410285829", -- LUT(4) = log10 (0.9991) = -0.00039104102858294304
--		x"0000390882623694", -- LUT(5) = log10 (0.99991) = -0.000039088262369485056
--		x"0000039086679261", -- LUT(6) = log10 (0.999991) = -0.0000039086679261613178
--		x"0000003908652096", -- LUT(7) = log10 (0.9999991) = -3.9086520960229735E-7
--		x"0000000390865051", -- LUT(8) = log10 (0.99999991) = -3.9086505130185422E-8
--		x"0000000039086503", -- LUT(9) = log10 (0.999999991) = -3.9086503547181931E-9
--		x"0000000003908650", -- LUT(10) = log10 (0.9999999991) = -3.9086503388881591E-10
--		x"0000000000390865", -- LUT(11) = log10 (0.99999999991) = -3.9086503373051557E-11
--		x"0000000000039086", -- LUT(12) = log10 (0.999999999991) = -3.9086503371468554E-12
--		x"0000000000003908", -- LUT(13) = log10 (0.9999999999991) = -3.9086503371310253E-13
--		x"0000000000000390", -- LUT(14) = log10 (0.99999999999991) = -3.9086503371294423E-14
--		x"0000000000000039"); -- LUT(15) = log10 (0.999999999999991) = -3.9086503371292840E-15

--
--signal lut_Log10ShP1: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"0457574905606751254099441934897693", -- LUT(1) = log10 (0.9) = -0.045757490560675125409944193489769382
--		x"0043648054024500846597442222467451", -- LUT(2) = log10 (0.99) = -0.0043648054024500846597442222467451399
--		x"0004345117740176913064656006955246", -- LUT(3) = log10 (0.999) = -0.00043451177401769130646560069552462442
--		x"0000434316198075103845560440238072", -- LUT(4) = log10 (0.9999) = -0.000043431619807510384556044023807226674
--		x"0000043429665339013793521486464083", -- LUT(5) = log10 (0.99999) = -0.0000043429665339013793521486464083130412
--		x"0000004342946990506375442129175357", -- LUT(6) = log10 (0.999999) = -4.3429469905063754421291753575839664E-7
--		x"0000000434294503617977370462101885", -- LUT(7) = log10 (0.9999999) = -4.3429450361797737046210188594163824E-8
--		x"0000000043429448407472425164387089", -- LUT(8) = log10 (0.99999999) = -4.3429448407472425164387089585426528E-9
--		x"0000000004342944821203990687475196", -- LUT(9) = log10 (0.999999999) = -4.3429448212039906874751966015182710E-10
--		x"0000000000434294481924966551747739", -- LUT(10) = log10 (0.9999999999) = -4.3429448192496655174773915857228094E-11
--		x"0000000000043429448190542330006065", -- LUT(11) = log10 (0.99999999999) = -4.3429448190542330006065965453759094E-12
--		x"0000000000004342944819034689748920", -- LUT(12) = log10 (0.999999999999) = -4.3429448190346897489208068959525795E-13
--		x"0000000000000434294481903273542375", -- LUT(13) = log10 (0.9999999999999) = -4.3429448190327354237522408295563591E-14
--		x"0000000000000043429448190325399912", -- LUT(14) = log10 (0.99999999999999) = -4.3429448190325399912353843519021982E-15
--		x"0000000000000004342944819032520447", -- LUT(15) = log10 (0.999999999999999) = -4.3429448190325204479836987054266367E-16
--		x"0000000000000000434294481903251849", -- LUT(16) = log10 (0.9999999999999999) = -4.3429448190325184936585301407919791E-17
--		x"0000000000000000043429448190325182", -- LUT(17) = log10 (0.99999999999999999) = -4.3429448190325182982260132843286424E-18
--		x"0000000000000000004342944819032518", -- LUT(18) = log10 (0.999999999999999999) = -4.3429448190325182786827615986823100E-19
--		x"0000000000000000000434294481903251", -- LUT(19) = log10 (0.9999999999999999999) = -4.3429448190325182767284364301176767E-20
--		x"0000000000000000000043429448190325", -- LUT(20) = log10 (0.99999999999999999999) = -4.3429448190325182765330039132612134E-21
--		x"0000000000000000000004342944819032", -- LUT(21) = log10 (0.999999999999999999999) = -4.3429448190325182765134606615755671E-22
--		x"0000000000000000000000434294481903", -- LUT(22) = log10 (0.9999999999999999999999) = -4.3429448190325182765115063364070024E-23
--		x"0000000000000000000000043429448190", -- LUT(23) = log10 (0.99999999999999999999999) = -4.3429448190325182765113109038901460E-24
--		x"0000000000000000000000004342944819", -- LUT(24) = log10 (0.999999999999999999999999) = -4.3429448190325182765112913606384603E-25
--		x"0000000000000000000000000434294481", -- LUT(25) = log10 (0.9999999999999999999999999) = -4.3429448190325182765112894063132918E-26
--		x"0000000000000000000000000043429448", -- LUT(26) = log10 (0.99999999999999999999999999) = -4.3429448190325182765112892108807749E-27
--		x"0000000000000000000000000004342944", -- LUT(27) = log10 (0.999999999999999999999999999) = -4.3429448190325182765112891913375232E-28
--		x"0000000000000000000000000000434294", -- LUT(28) = log10 (0.9999999999999999999999999999) = -4.3429448190325182765112891893831981E-29
--		x"0000000000000000000000000000043429", -- LUT(29) = log10 (0.99999999999999999999999999999) = -4.3429448190325182765112891891877655E-30
--		x"0000000000000000000000000000004342", -- LUT(30) = log10 (0.999999999999999999999999999999) = -4.3429448190325182765112891891682223E-31
--		x"0000000000000000000000000000000434", -- LUT(31) = log10 (0.9999999999999999999999999999999) = -4.3429448190325182765112891891662680E-32
--		x"0000000000000000000000000000000043", -- LUT(32) = log10 (0.99999999999999999999999999999999) = -4.3429448190325182765112891891660725E-33
--		x"0000000000000000000000000000000004"); -- LUT(33) = log10 (0.999999999999999999999999999999999) = -4.3429448190325182765112891891660530E-34
--
--signal lut_Log10ShP2: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"0969100130080564143587833158265209", -- LUT(1) = log10 (0.8) = -0.096910013008056414358783315826520920
--		x"0087739243075051433618285880902345", -- LUT(2) = log10 (0.98) = -0.0087739243075051433618285880902345863
--		x"0008694587126288906203560692421185", -- LUT(3) = log10 (0.998) = -0.00086945871262889062035606924211850592
--		x"0000868675834285807945676917580550", -- LUT(4) = log10 (0.9998) = -0.000086867583428580794567691758055002046
--		x"0000086859764981195531938540093755", -- LUT(5) = log10 (0.99998) = -0.0000086859764981195531938540093755639715
--		x"0000008685898323966255821615025187", -- LUT(6) = log10 (0.999998) = -8.6858983239662558216150251873377498E-7
--		x"0000000868589050665411617140544632", -- LUT(7) = log10 (0.9999998) = -8.6858905066541161714054463297995950E-8
--		x"0000000086858897249239340917915796", -- LUT(8) = log10 (0.99999998) = -8.6858897249239340917915796890089799E-9
--		x"0000000008685889646750926202668801", -- LUT(9) = log10 (0.999999998) = -8.6858896467509262026688011328131747E-10
--		x"0000000000868588963893362551694489", -- LUT(10) = log10 (0.9999999998) = -8.6858896389336255169448938954925984E-11
--		x"0000000000086858896381518954494043", -- LUT(11) = log10 (0.99999999998) = -8.6858896381518954494043868624807535E-12
--		x"0000000000008685889638073722442660", -- LUT(12) = log10 (0.999999999998) = -8.6858896380737224426606549960713083E-13
--		x"0000000000000868588963806590514198", -- LUT(13) = log10 (0.9999999999998) = -8.6858896380659051419863849977992657E-14
--		x"0000000000000086858896380651234119", -- LUT(14) = log10 (0.99999999999998) = -8.6858896380651234119189590298557505E-15
--		x"0000000000000008685889638065045238", -- LUT(15) = log10 (0.999999999999998) = -8.6858896380650452389122164433802359E-16
--		x"0000000000000000868588963806503742", -- LUT(16) = log10 (0.9999999999999998) = -8.6858896380650374216115421848358728E-17
--		x"0000000000000000086858896380650366", -- LUT(17) = log10 (0.99999999999999998) = -8.6858896380650366398814747589824683E-18
--		x"0000000000000000008685889638065036", -- LUT(18) = log10 (0.999999999999999998) = -8.6858896380650365617084680163971382E-19
--		x"0000000000000000000868588963806503", -- LUT(19) = log10 (0.9999999999999999998) = -8.6858896380650365538911673421386053E-20
--		x"0000000000000000000086858896380650", -- LUT(20) = log10 (0.99999999999999999998) = -8.6858896380650365531094372747127520E-21
--		x"0000000000000000000008685889638065", -- LUT(21) = log10 (0.999999999999999999998) = -8.6858896380650365530312642679701667E-22
--		x"0000000000000000000000868588963806", -- LUT(22) = log10 (0.9999999999999999999998) = -8.6858896380650365530234469672959081E-23
--		x"0000000000000000000000086858896380", -- LUT(23) = log10 (0.99999999999999999999998) = -8.6858896380650365530226652372284823E-24
--		x"0000000000000000000000008685889638", -- LUT(24) = log10 (0.999999999999999999999998) = -8.6858896380650365530225870642217397E-25
--		x"0000000000000000000000000868588963", -- LUT(25) = log10 (0.9999999999999999999999998) = -8.6858896380650365530225792469210655E-26
--		x"0000000000000000000000000086858896", -- LUT(26) = log10 (0.99999999999999999999999998) = -8.6858896380650365530225784651909980E-27
--		x"0000000000000000000000000008685889", -- LUT(27) = log10 (0.999999999999999999999999998) = -8.6858896380650365530225783870179913E-28
--		x"0000000000000000000000000000868588", -- LUT(28) = log10 (0.9999999999999999999999999998) = -8.6858896380650365530225783792006906E-29
--		x"0000000000000000000000000000086858", -- LUT(29) = log10 (0.99999999999999999999999999998) = -8.6858896380650365530225783784189605E-30
--		x"0000000000000000000000000000008685", -- LUT(30) = log10 (0.999999999999999999999999999998) = -8.6858896380650365530225783783407875E-31
--		x"0000000000000000000000000000000868", -- LUT(31) = log10 (0.9999999999999999999999999999998) = -8.6858896380650365530225783783329702E-32
--		x"0000000000000000000000000000000086", -- LUT(32) = log10 (0.99999999999999999999999999999998) = -8.6858896380650365530225783783321885E-33
--		x"0000000000000000000000000000000008"); -- LUT(33) = log10 (0.999999999999999999999999999999998) = -8.6858896380650365530225783783321103E-34
--
--signal lut_Log10ShP3: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"1549019599857431692877837414073638", -- LUT(1) = log10 (0.7) = -0.15490195998574316928778374140736381
--		x"0132282657337551482156381883344225", -- LUT(2) = log10 (0.97) = -0.013228265733755148215638188334422551
--		x"0013048416883442801186282971867276", -- LUT(3) = log10 (0.997) = -0.0013048416883442801186282971867276073
--		x"0001303078917321911892026020669822", -- LUT(4) = log10 (0.9997) = -0.00013030789173219118920260206698228363
--		x"0000130290298935231495767288863830", -- LUT(5) = log10 (0.99997) = -0.000013029029893523149576728886383053175
--		x"0000013028854000388327067182248185", -- LUT(6) = log10 (0.999997) = -0.0000013028854000388327067182248185842475
--		x"0000001302883641142311425928874957", -- LUT(7) = log10 (0.9999997) = -1.3028836411423114259288749577915299E-7
--		x"0000000130288346525300755946476150", -- LUT(8) = log10 (0.99999997) = -1.3028834652530075594647615084407311E-8
--		x"0000000013028834476640806554266703", -- LUT(9) = log10 (0.999999997) = -1.3028834476640806554266703271036251E-9
--		x"0000000001302883445905187999848936", -- LUT(10) = log10 (0.9999999997) = -1.3028834459051879998489365825729104E-10
--		x"0000000000130288344572929873463942", -- LUT(11) = log10 (0.99999999997) = -1.3028834457292987346394239540278378E-11
--		x"0000000000013028834457117098081219", -- LUT(12) = log10 (0.999999999997) = -1.3028834457117098081219552986245825E-12
--		x"0000000000001302883445709950915470", -- LUT(13) = log10 (0.9999999999997) = -1.3028834457099509154702432591587616E-13
--		x"0000000000000130288344570977502620", -- LUT(14) = log10 (0.99999999999997) = -1.3028834457097750262050724034729246E-14
--		x"0000000000000013028834457097574372", -- LUT(15) = log10 (0.999999999999997) = -1.3028834457097574372785553213869483E-15
--		x"0000000000000001302883445709755678", -- LUT(16) = log10 (0.9999999999999997) = -1.3028834457097556783859036132131768E-16
--		x"0000000000000000130288344570975550", -- LUT(17) = log10 (0.99999999999999997) = -1.3028834457097555024966384423961479E-17
--		x"0000000000000000013028834457097554", -- LUT(18) = log10 (0.999999999999999997) = -1.3028834457097554849077119253144485E-18
--		x"0000000000000000001302883445709755", -- LUT(19) = log10 (0.9999999999999999997) = -1.3028834457097554831488192736062786E-19
--		x"0000000000000000000130288344570975", -- LUT(20) = log10 (0.99999999999999999997) = -1.3028834457097554829729300084354616E-20
--		x"0000000000000000000013028834457097", -- LUT(21) = log10 (0.999999999999999999997) = -1.3028834457097554829553410819183799E-21
--		x"0000000000000000000001302883445709", -- LUT(22) = log10 (0.9999999999999999999997) = -1.3028834457097554829535821892666717E-22
--		x"0000000000000000000000130288344570", -- LUT(23) = log10 (0.99999999999999999999997) = -1.3028834457097554829534063000015009E-23
--		x"0000000000000000000000013028834457", -- LUT(24) = log10 (0.999999999999999999999997) = -1.3028834457097554829533887110749838E-24
--		x"0000000000000000000000001302883445", -- LUT(25) = log10 (0.9999999999999999999999997) = -1.3028834457097554829533869521823321E-25
--		x"0000000000000000000000000130288344", -- LUT(26) = log10 (0.99999999999999999999999997) = -1.3028834457097554829533867762930669E-26
--		x"0000000000000000000000000013028834", -- LUT(27) = log10 (0.999999999999999999999999997) = -1.3028834457097554829533867587041404E-27
--		x"0000000000000000000000000001302883", -- LUT(28) = log10 (0.9999999999999999999999999997) = -1.3028834457097554829533867569452478E-28
--		x"0000000000000000000000000000130288", -- LUT(29) = log10 (0.99999999999999999999999999997) = -1.3028834457097554829533867567693585E-29
--		x"0000000000000000000000000000013028", -- LUT(30) = log10 (0.999999999999999999999999999997) = -1.3028834457097554829533867567517696E-30
--		x"0000000000000000000000000000001302", -- LUT(31) = log10 (0.9999999999999999999999999999997) = -1.3028834457097554829533867567500107E-31
--		x"0000000000000000000000000000000130", -- LUT(32) = log10 (0.99999999999999999999999999999997) = -1.3028834457097554829533867567498348E-32
--		x"0000000000000000000000000000000013"); -- LUT(33) = log10 (0.999999999999999999999999999999997) = -1.3028834457097554829533867567498172E-33
--
--signal lut_Log10ShP4: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"2218487496163563674912332020203916", -- LUT(1) = log10 (0.6) = -0.22184874961635636749123320202039166
--		x"0177287669604315866362776231224195", -- LUT(2) = log10 (0.96) = -0.017728766960431586636277623122419557
--		x"0017406615763012684447339552686373", -- LUT(3) = log10 (0.996) = -0.0017406615763012684447339552686373903
--		x"0001737525455875823128918957822892", -- LUT(4) = log10 (0.9996) = -0.00017375254558758231289189578228922029
--		x"0000173721267209808226121397155421", -- LUT(5) = log10 (0.99996) = -0.000017372126720980822612139715542103355
--		x"0000017371814019781275133613420426", -- LUT(6) = log10 (0.999996) = -0.0000017371814019781275133613420426354859
--		x"0000001737178275048685482723245346", -- LUT(7) = log10 (0.9999996) = -1.7371782750486854827232453460289498E-7
--		x"0000000173717796235656678935958440", -- LUT(8) = log10 (0.99999996) = -1.7371779623565667893595844095416974E-8
--		x"0000000017371779310873631750954792", -- LUT(9) = log10 (0.999999996) = -1.7371779310873631750954792719396709E-9
--		x"0000000001737177927960442896219766", -- LUT(10) = log10 (0.9999999996) = -1.7371779279604428962197666272878120E-10
--		x"0000000000173717792764775086915770", -- LUT(11) = log10 (0.99999999996) = -1.7371779276477508691577023167732654E-11
--		x"0000000000017371779276164816664597", -- LUT(12) = log10 (0.999999999996) = -1.7371779276164816664597509552365767E-12
--		x"0000000000001737177927613354746190", -- LUT(13) = log10 (0.9999999999996) = -1.7371779276133547461900383697780307E-13
--		x"0000000000000173717792761304205416", -- LUT(14) = log10 (0.99999999999996) = -1.7371779276130420541630679367391273E-14
--		x"0000000000000017371779276130107849", -- LUT(15) = log10 (0.999999999999996) = -1.7371779276130107849603709016903065E-15
--		x"0000000000000001737177927613007658", -- LUT(16) = log10 (0.9999999999999996) = -1.7371779276130076580401011982679751E-16
--		x"0000000000000000173717792761300734", -- LUT(17) = log10 (0.99999999999999996) = -1.7371779276130073453480742279265675E-17
--		x"0000000000000000017371779276130073", -- LUT(18) = log10 (0.999999999999999996) = -1.7371779276130073140788715308924350E-18
--		x"0000000000000000001737177927613007", -- LUT(19) = log10 (0.9999999999999999996) = -1.7371779276130073109519512611890218E-19
--		x"0000000000000000000173717792761300", -- LUT(20) = log10 (0.99999999999999999996) = -1.7371779276130073106392592342186805E-20
--		x"0000000000000000000017371779276130", -- LUT(21) = log10 (0.999999999999999999996) = -1.7371779276130073106079900315216463E-21
--		x"0000000000000000000001737177927613", -- LUT(22) = log10 (0.9999999999999999999996) = -1.7371779276130073106048631112519429E-22
--		x"0000000000000000000000173717792761", -- LUT(23) = log10 (0.99999999999999999999996) = -1.7371779276130073106045504192249726E-23
--		x"0000000000000000000000017371779276", -- LUT(24) = log10 (0.999999999999999999999996) = -1.7371779276130073106045191500222756E-24
--		x"0000000000000000000000001737177927", -- LUT(25) = log10 (0.9999999999999999999999996) = -1.7371779276130073106045160231020059E-25
--		x"0000000000000000000000000173717792", -- LUT(26) = log10 (0.99999999999999999999999996) = -1.7371779276130073106045157104099789E-26
--		x"0000000000000000000000000017371779", -- LUT(27) = log10 (0.999999999999999999999999996) = -1.7371779276130073106045156791407762E-27
--		x"0000000000000000000000000001737177", -- LUT(28) = log10 (0.9999999999999999999999999996) = -1.7371779276130073106045156760138559E-28
--		x"0000000000000000000000000000173717", -- LUT(29) = log10 (0.99999999999999999999999999996) = -1.7371779276130073106045156757011639E-29
--		x"0000000000000000000000000000017371", -- LUT(30) = log10 (0.999999999999999999999999999996) = -1.7371779276130073106045156756698947E-30
--		x"0000000000000000000000000000001737", -- LUT(31) = log10 (0.9999999999999999999999999999996) = -1.7371779276130073106045156756667678E-31
--		x"0000000000000000000000000000000173", -- LUT(32) = log10 (0.99999999999999999999999999999996) = -1.7371779276130073106045156756664551E-32
--		x"0000000000000000000000000000000017"); -- LUT(33) = log10 (0.999999999999999999999999999999996) = -1.7371779276130073106045156756664238E-33
--
--signal lut_Log10ShP5: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"3010299956639811952137388947244930", -- LUT(1) = log10 (0.5) = -0.30102999566398119521373889472449303
--		x"0222763947111522336774054189675637", -- LUT(2) = log10 (0.95) = -0.022276394711152233677405418967563709
--		x"0021769192542745451137171103046901", -- LUT(3) = log10 (0.995) = -0.0021769192542745451137171103046901853
--		x"0002172015458642557996912240036058", -- LUT(4) = log10 (0.9995) = -0.00021720154586425579969122400360587672
--		x"0000217152669813612524722490126493", -- LUT(5) = log10 (0.99995) = -0.000021715266981361252472249012649395659
--		x"0000021714778382153786001749099590", -- LUT(6) = log10 (0.999995) = -0.0000021714778382153786001749099590785766
--		x"0000002171472952384542473422414053", -- LUT(7) = log10 (0.9999995) = -2.1714729523845424734224140533631616E-7
--		x"0000000217147246380307118572253217", -- LUT(8) = log10 (0.99999995) = -2.1714724638030711857225321730389339E-8
--		x"0000000021714724149449401801418959", -- LUT(9) = log10 (0.999999995) = -2.1714724149449401801418959207161428E-9
--		x"0000000002171472410059127240815665", -- LUT(10) = log10 (0.9999999995) = -2.1714724100591272408156654133411500E-10
--		x"0000000000217147240957054594849536", -- LUT(11) = log10 (0.99999999995) = -2.1714724095705459484953606333807479E-11
--		x"0000000000021714724095216878192794", -- LUT(12) = log10 (0.999999999995) = -2.1714724095216878192794533380320772E-12
--		x"0000000000002171472409516802006358", -- LUT(13) = log10 (0.9999999999995) = -2.1714724095168020063580238403236234E-13
--		x"0000000000000217147240951631342506", -- LUT(14) = log10 (0.99999999999995) = -2.1714724095163134250658825028710421E-14
--		x"0000000000000021714724095162645669", -- LUT(15) = log10 (0.999999999999995) = -2.1714724095162645669366683852489667E-15
--		x"0000000000000002171472409516259681", -- LUT(16) = log10 (0.9999999999999995) = -2.1714724095162596811237469736479909E-16
--		x"0000000000000000217147240951625919", -- LUT(17) = log10 (0.99999999999999995) = -2.1714724095162591925424548324895057E-17
--		x"0000000000000000021714724095162591", -- LUT(18) = log10 (0.999999999999999995) = -2.1714724095162591436843256183736733E-18
--		x"0000000000000000002171472409516259", -- LUT(19) = log10 (0.9999999999999999995) = -2.1714724095162591387985126969620902E-19
--		x"0000000000000000000217147240951625", -- LUT(20) = log10 (0.99999999999999999995) = -2.1714724095162591383099314048209319E-20
--		x"0000000000000000000021714724095162", -- LUT(21) = log10 (0.999999999999999999995) = -2.1714724095162591382610732756068161E-21
--		x"0000000000000000000002171472409516", -- LUT(22) = log10 (0.9999999999999999999995) = -2.1714724095162591382561874626854045E-22
--		x"0000000000000000000000217147240951", -- LUT(23) = log10 (0.99999999999999999999995) = -2.1714724095162591382556988813932633E-23
--		x"0000000000000000000000021714724095", -- LUT(24) = log10 (0.999999999999999999999995) = -2.1714724095162591382556500232640492E-24
--		x"0000000000000000000000002171472409", -- LUT(25) = log10 (0.9999999999999999999999995) = -2.1714724095162591382556451374511278E-25
--		x"0000000000000000000000000217147240", -- LUT(26) = log10 (0.99999999999999999999999995) = -2.1714724095162591382556446488698356E-26
--		x"0000000000000000000000000021714724", -- LUT(27) = log10 (0.999999999999999999999999995) = -2.1714724095162591382556446000117064E-27
--		x"0000000000000000000000000002171472", -- LUT(28) = log10 (0.9999999999999999999999999995) = -2.1714724095162591382556445951258935E-28
--		x"0000000000000000000000000000217147", -- LUT(29) = log10 (0.99999999999999999999999999995) = -2.1714724095162591382556445946373122E-29
--		x"0000000000000000000000000000021714", -- LUT(30) = log10 (0.999999999999999999999999999995) = -2.1714724095162591382556445945884541E-30
--		x"0000000000000000000000000000002171", -- LUT(31) = log10 (0.9999999999999999999999999999995) = -2.1714724095162591382556445945835683E-31
--		x"0000000000000000000000000000000217", -- LUT(32) = log10 (0.99999999999999999999999999999995) = -2.1714724095162591382556445945830797E-32
--		x"0000000000000000000000000000000021"); -- LUT(33) = log10 (0.999999999999999999999999999999995) = -2.1714724095162591382556445945830308E-33
--
--signal lut_Log10ShP6: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"3979400086720376095725222105510139", -- LUT(1) = log10 (0.4) = -0.39794000867203760957252221055101395
--		x"0268721464003013403720417058263063", -- LUT(2) = log10 (0.94) = -0.026872146400301340372041705826306333
--		x"0026136156026866879812154116474416", -- LUT(3) = log10 (0.994) = -0.0026136156026866879812154116474416445
--		x"0002606548934319742776940456484595", -- LUT(4) = log10 (0.9994) = -0.00026065489343197427769404564845954106
--		x"0000260584506755331453910578603670", -- LUT(5) = log10 (0.99994) = -0.000026058450675533145391057860367025435
--		x"0000026057747087514545678487929202", -- LUT(6) = log10 (0.999994) = -0.0000026057747087514545678487929202199916
--		x"0000002605767673149891083927745106", -- LUT(7) = log10 (0.9999994) = -2.6057676731498910839277451065257585E-7
--		x"0000000260576696959252083541251290", -- LUT(8) = log10 (0.99999994) = -2.6057669695925208354125129055348858E-8
--		x"0000000026057668992368116714345092", -- LUT(9) = log10 (0.999999994) = -2.6057668992368116714345092489654954E-9
--		x"0000000002605766892201241033645318", -- LUT(10) = log10 (0.9999999994) = -2.6057668922012410336453188303827153E-10
--		x"0000000000260576689149768397265248", -- LUT(11) = log10 (0.99999999994) = -2.6057668914976839726524857627466778E-11
--		x"0000000000026057668914273282665810", -- LUT(12) = log10 (0.999999999994) = -2.6057668914273282665810633156000480E-12
--		x"0000000000002605766891420292695974", -- LUT(13) = log10 (0.9999999999994) = -2.6057668914202926959741996794814295E-13
--		x"0000000000000260576689141958913891", -- LUT(14) = log10 (0.99999999999994) = -2.6057668914195891389135161019555280E-14
--		x"0000000000000026057668914195187832", -- LUT(15) = log10 (0.999999999999994) = -2.6057668914195187832074477720637974E-15
--		x"0000000000000002605766891419511747", -- LUT(16) = log10 (0.9999999999999994) = -2.6057668914195117476368409393532330E-16
--		x"0000000000000000260576689141951104", -- LUT(17) = log10 (0.99999999999999994) = -2.6057668914195110440797802560849626E-17
--		x"0000000000000000026057668914195109", -- LUT(18) = log10 (0.999999999999999994) = -2.6057668914195109737240741877581634E-18
--		x"0000000000000000002605766891419510", -- LUT(19) = log10 (0.9999999999999999994) = -2.6057668914195109666885035809254838E-19
--		x"0000000000000000000260576689141951", -- LUT(20) = log10 (0.99999999999999999994) = -2.6057668914195109659849465202422158E-20
--		x"0000000000000000000026057668914195", -- LUT(21) = log10 (0.999999999999999999994) = -2.6057668914195109659145908141738890E-21
--		x"0000000000000000000002605766891419", -- LUT(22) = log10 (0.9999999999999999999994) = -2.6057668914195109659075552435670563E-22
--		x"0000000000000000000000260576689141", -- LUT(23) = log10 (0.99999999999999999999994) = -2.6057668914195109659068516865063731E-23
--		x"0000000000000000000000026057668914", -- LUT(24) = log10 (0.999999999999999999999994) = -2.6057668914195109659067813308003048E-24
--		x"0000000000000000000000002605766891", -- LUT(25) = log10 (0.9999999999999999999999994) = -2.6057668914195109659067742952296979E-25
--		x"0000000000000000000000000260576689", -- LUT(26) = log10 (0.99999999999999999999999994) = -2.6057668914195109659067735916726372E-26
--		x"0000000000000000000000000026057668", -- LUT(27) = log10 (0.999999999999999999999999994) = -2.6057668914195109659067735213169312E-27
--		x"0000000000000000000000000002605766", -- LUT(28) = log10 (0.9999999999999999999999999994) = -2.6057668914195109659067735142813606E-28
--		x"0000000000000000000000000000260576", -- LUT(29) = log10 (0.99999999999999999999999999994) = -2.6057668914195109659067735135778035E-29
--		x"0000000000000000000000000000026057", -- LUT(30) = log10 (0.999999999999999999999999999994) = -2.6057668914195109659067735135074478E-30
--		x"0000000000000000000000000000002605", -- LUT(31) = log10 (0.9999999999999999999999999999994) = -2.6057668914195109659067735135004122E-31
--		x"0000000000000000000000000000000260", -- LUT(32) = log10 (0.99999999999999999999999999999994) = -2.6057668914195109659067735134997087E-32
--		x"0000000000000000000000000000000026"); -- LUT(33) = log10 (0.999999999999999999999999999999994) = -2.6057668914195109659067735134996383E-33
--
--signal lut_Log10ShP7: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"5228787452803375627049720967448846", -- LUT(1) = log10 (0.3) = -0.52287874528033756270497209674488469
--		x"0315170514460648830382679966264689", -- LUT(2) = log10 (0.93) = -0.031517051446064883038267996626468968
--		x"0030507515046188240968314894040280", -- LUT(3) = log10 (0.993) = -0.0030507515046188240968314894040280557
--		x"0003041125891607614734971455976653", -- LUT(4) = log10 (0.9993) = -0.00030411258916076147349714559766534881
--		x"0000304016778043652336654484495304", -- LUT(5) = log10 (0.99993) = -0.000030401677804365233665448449530405305
--		x"0000030400720135872240196786742857", -- LUT(6) = log10 (0.999993) = -0.0000030400720135872240196786742857836769
--		x"0000003040062437344740000143208304", -- LUT(7) = log10 (0.9999993) = -3.0400624373447400001432083043512939E-7
--		x"0000000304006147972491582528843731", -- LUT(8) = log10 (0.99999993) = -3.0400614797249158252884373193994110E-8
--		x"0000000030400613839629776498419082", -- LUT(9) = log10 (0.999999993) = -3.0400613839629776498419082348259506E-9
--		x"0000000003040061374386784274717412", -- LUT(10) = log10 (0.9999999993) = -3.0400613743867842747174127680649046E-10
--		x"0000000000304006137342916494162916", -- LUT(11) = log10 (0.99999999993) = -3.0400613734291649416291645637674500E-11
--		x"0000000000030400613733334030083645", -- LUT(12) = log10 (0.999999999993) = -3.0400613733334030083645817565294528E-12
--		x"0000000000003040061373323826815038", -- LUT(13) = log10 (0.9999999999993) = -3.0400613733238268150385658959373385E-13
--		x"0000000000000304006137332286919570", -- LUT(14) = log10 (0.99999999999993) = -3.0400613733228691957059687340794437E-14
--		x"0000000000000030400613733227734337", -- LUT(15) = log10 (0.999999999999993) = -3.0400613733227734337727090621356674E-15
--		x"0000000000000003040061373322763857", -- LUT(16) = log10 (0.9999999999999993) = -3.0400613733227638575793830953837099E-16
--		x"0000000000000000304006137332276289", -- LUT(17) = log10 (0.99999999999999993) = -3.0400613733227628999600504987129383E-17
--		x"0000000000000000030400613733227628", -- LUT(18) = log10 (0.999999999999999993) = -3.0400613733227628041981172390459054E-18
--		x"0000000000000000003040061373322762", -- LUT(19) = log10 (0.9999999999999999993) = -3.0400613733227627946219239130792026E-19
--		x"0000000000000000000304006137332276", -- LUT(20) = log10 (0.99999999999999999993) = -3.0400613733227627936643045804825323E-20
--		x"0000000000000000000030400613733227", -- LUT(21) = log10 (0.999999999999999999993) = -3.0400613733227627935685426472228652E-21
--		x"0000000000000000000003040061373322", -- LUT(22) = log10 (0.9999999999999999999993) = -3.0400613733227627935589664538968985E-22
--		x"0000000000000000000000304006137332", -- LUT(23) = log10 (0.99999999999999999999993) = -3.0400613733227627935580088345643019E-23
--		x"0000000000000000000000030400613733", -- LUT(24) = log10 (0.999999999999999999999993) = -3.0400613733227627935579130726310422E-24
--		x"0000000000000000000000003040061373", -- LUT(25) = log10 (0.9999999999999999999999993) = -3.0400613733227627935579034964377162E-25
--		x"0000000000000000000000000304006137", -- LUT(26) = log10 (0.99999999999999999999999993) = -3.0400613733227627935579025388183836E-26
--		x"0000000000000000000000000030400613", -- LUT(27) = log10 (0.999999999999999999999999993) = -3.0400613733227627935579024430564504E-27
--		x"0000000000000000000000000003040061", -- LUT(28) = log10 (0.9999999999999999999999999993) = -3.0400613733227627935579024334802571E-28
--		x"0000000000000000000000000000304006", -- LUT(29) = log10 (0.99999999999999999999999999993) = -3.0400613733227627935579024325226377E-29
--		x"0000000000000000000000000000030400", -- LUT(30) = log10 (0.999999999999999999999999999993) = -3.0400613733227627935579024324268758E-30
--		x"0000000000000000000000000000003040", -- LUT(31) = log10 (0.9999999999999999999999999999993) = -3.0400613733227627935579024324172996E-31
--		x"0000000000000000000000000000000304", -- LUT(32) = log10 (0.99999999999999999999999999999993) = -3.0400613733227627935579024324163420E-32
--		x"0000000000000000000000000000000030"); -- LUT(33) = log10 (0.999999999999999999999999999999993) = -3.0400613733227627935579024324162462E-33
--
--signal lut_Log10ShP8: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"6989700043360188047862611052755069", -- LUT(1) = log10 (0.2) = -0.69897000433601880478626110527550697
--		x"0362121726544447307047450982998243", -- LUT(2) = log10 (0.92) = -0.036212172654444730704745098299824397
--		x"0034883278458213442646014262591191", -- LUT(3) = log10 (0.992) = -0.0034883278458213442646014262591191439
--		x"0003475746339209023167184248040235", -- LUT(4) = log10 (0.9992) = -0.00034757463392090231671842480402357271
--		x"0000347449483687262756562266725871", -- LUT(5) = log10 (0.99992) = -0.000034744948368726275656226672587143454
--		x"0000034743697527235555615660668462", -- LUT(6) = log10 (0.999992) = -0.0000034743697527235555615660668462652569
--		x"0000003474357244969097907975379218", -- LUT(7) = log10 (0.9999992) = -3.4743572449690979079753792188195904E-7
--		x"0000000347435599420025624220921873", -- LUT(8) = log10 (0.99999992) = -3.4743559942002562422092187327698841E-8
--		x"0000000034743558691234381162326818", -- LUT(9) = log10 (0.999999992) = -3.4743558691234381162326818590414970E-9
--		x"0000000003474355856615756964040633", -- LUT(10) = log10 (0.9999999992) = -3.4743558566157569640406331160427205E-10
--		x"0000000000347435585536498885542548", -- LUT(11) = log10 (0.99999999992) = -3.4743558553649888554254838953394621E-11
--		x"0000000000034743558552399120446300", -- LUT(12) = log10 (0.999999999992) = -3.4743558552399120446300095294092554E-12
--		x"0000000000003474355855227404363551", -- LUT(13) = log10 (0.9999999999992) = -3.4743558552274043635511224983772401E-13
--		x"0000000000000347435585522615359544", -- LUT(14) = log10 (0.99999999999992) = -3.4743558552261535954432403993296482E-14
--		x"0000000000000034743558552260285186", -- LUT(15) = log10 (0.999999999999992) = -3.4743558552260285186324522554654451E-15
--		x"0000000000000003474355855226016010", -- LUT(16) = log10 (0.9999999999999992) = -3.4743558552260160109513734417394303E-16
--		x"0000000000000000347435585522601476", -- LUT(17) = log10 (0.99999999999999992) = -3.4743558552260147601832655603734329E-17
--		x"0000000000000000034743558552260146", -- LUT(18) = log10 (0.999999999999999992) = -3.4743558552260146351064547722368992E-18
--		x"0000000000000000003474355855226014", -- LUT(19) = log10 (0.9999999999999999992) = -3.4743558552260146225987736934232465E-19
--		x"0000000000000000000347435585522601", -- LUT(20) = log10 (0.99999999999999999992) = -3.4743558552260146213480055855418812E-20
--		x"0000000000000000000034743558552260", -- LUT(21) = log10 (0.999999999999999999992) = -3.4743558552260146212229287747537447E-21
--		x"0000000000000000000003474355855226", -- LUT(22) = log10 (0.9999999999999999999992) = -3.4743558552260146212104210936749311E-22
--		x"0000000000000000000000347435585522", -- LUT(23) = log10 (0.99999999999999999999992) = -3.4743558552260146212091703255670497E-23
--		x"0000000000000000000000034743558552", -- LUT(24) = log10 (0.999999999999999999999992) = -3.4743558552260146212090452487562616E-24
--		x"0000000000000000000000003474355855", -- LUT(25) = log10 (0.9999999999999999999999992) = -3.4743558552260146212090327410751827E-25
--		x"0000000000000000000000000347435585", -- LUT(26) = log10 (0.99999999999999999999999992) = -3.4743558552260146212090314903070749E-26
--		x"0000000000000000000000000034743558", -- LUT(27) = log10 (0.999999999999999999999999992) = -3.4743558552260146212090313652302641E-27
--		x"0000000000000000000000000003474355", -- LUT(28) = log10 (0.9999999999999999999999999992) = -3.4743558552260146212090313527225830E-28
--		x"0000000000000000000000000000347435", -- LUT(29) = log10 (0.99999999999999999999999999992) = -3.4743558552260146212090313514718149E-29
--		x"0000000000000000000000000000034743", -- LUT(30) = log10 (0.999999999999999999999999999992) = -3.4743558552260146212090313513467381E-30
--		x"0000000000000000000000000000003474", -- LUT(31) = log10 (0.9999999999999999999999999999992) = -3.4743558552260146212090313513342304E-31
--		x"0000000000000000000000000000000347", -- LUT(32) = log10 (0.99999999999999999999999999999992) = -3.4743558552260146212090313513329796E-32
--		x"0000000000000000000000000000000034"); -- LUT(33) = log10 (0.999999999999999999999999999999992) = -3.4743558552260146212090313513328546E-33
--
--signal lut_Log10ShP9: mlut_LogShP := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"0000000000000000000000000000000000", -- LUT(1) = log10 (0.1) = -1
--		x"0409586076789064000812785834650353", -- LUT(2) = log10 (0.91) = -0.040958607678906400081278583465035376
--		x"0039263455147246716355656211845791", -- LUT(3) = log10 (0.991) = -0.0039263455147246716355656211845791359
--		x"0003910410285829430445669937541831", -- LUT(4) = log10 (0.9991) = -0.00039104102858294304456699375418312618
--		x"0000390882623694850557891647691700", -- LUT(5) = log10 (0.99991) = -0.000039088262369485055789164769170025271
--		x"0000039086679261613178020183232463", -- LUT(6) = log10 (0.999991) = -0.0000039086679261613178020183232463383566
--		x"0000003908652096022973493333439196", -- LUT(7) = log10 (0.9999991) = -3.9086520960229734933334391960980503E-7
--		x"0000000390865051301854217303377306", -- LUT(8) = log10 (0.99999991) = -3.9086505130185421730337730695513009E-8
--		x"0000000039086503547181930714754191", -- LUT(9) = log10 (0.999999991) = -3.9086503547181930714754191049618901E-9
--		x"0000000003908650338888159101623665", -- LUT(10) = log10 (0.9999999991) = -3.9086503388881591016236657639737713E-10
--		x"0000000000390865033730515571404153", -- LUT(11) = log10 (0.99999999991) = -3.9086503373051557140415306163591143E-11
--		x"0000000000039086503371468553753773", -- LUT(12) = log10 (0.999999999991) = -3.9086503371468553753773475028284197E-12
--		x"0000000000003908650337131025341511", -- LUT(13) = log10 (0.9999999999991) = -3.9086503371310253415118694954870238E-13
--		x"0000000000000390865033712944233812", -- LUT(14) = log10 (0.99999999999991) = -3.9086503371294423381253310977930004E-14
--		x"0000000000000039086503371292840377", -- LUT(15) = log10 (0.999999999999991) = -3.9086503371292840377866773520539992E-15
--		x"0000000000000003908650337129268207", -- LUT(16) = log10 (0.9999999999999991) = -3.9086503371292682077528119784204031E-16
--		x"0000000000000000390865033712926662", -- LUT(17) = log10 (0.99999999999999991) = -3.9086503371292666247494254410664465E-17
--		x"0000000000000000039086503371292664", -- LUT(18) = log10 (0.999999999999999991) = -3.9086503371292664664490867873311449E-18
--		x"0000000000000000003908650337129266", -- LUT(19) = log10 (0.9999999999999999991) = -3.9086503371292664506190529219576156E-19
--		x"0000000000000000000390865033712926", -- LUT(20) = log10 (0.99999999999999999991) = -3.9086503371292664490360495354202627E-20
--		x"0000000000000000000039086503371292", -- LUT(21) = log10 (0.999999999999999999991) = -3.9086503371292664488777491967665274E-21
--		x"0000000000000000000003908650337129", -- LUT(22) = log10 (0.9999999999999999999991) = -3.9086503371292664488619191629011539E-22
--		x"0000000000000000000000390865033712", -- LUT(23) = log10 (0.99999999999999999999991) = -3.9086503371292664488603361595146166E-23
--		x"0000000000000000000000039086503371", -- LUT(24) = log10 (0.999999999999999999999991) = -3.9086503371292664488601778591759628E-24
--		x"0000000000000000000000003908650337", -- LUT(25) = log10 (0.9999999999999999999999991) = -3.9086503371292664488601620291420974E-25
--		x"0000000000000000000000000390865033", -- LUT(26) = log10 (0.99999999999999999999999991) = -3.9086503371292664488601604461387109E-26
--		x"0000000000000000000000000039086503", -- LUT(27) = log10 (0.999999999999999999999999991) = -3.9086503371292664488601602878383723E-27
--		x"0000000000000000000000000003908650", -- LUT(28) = log10 (0.9999999999999999999999999991) = -3.9086503371292664488601602720083384E-28
--		x"0000000000000000000000000000390865", -- LUT(29) = log10 (0.99999999999999999999999999991) = -3.9086503371292664488601602704253350E-29
--		x"0000000000000000000000000000039086", -- LUT(30) = log10 (0.999999999999999999999999999991) = -3.9086503371292664488601602702670347E-30
--		x"0000000000000000000000000000003908", -- LUT(31) = log10 (0.9999999999999999999999999999991) = -3.9086503371292664488601602702512046E-31
--		x"0000000000000000000000000000000390", -- LUT(32) = log10 (0.99999999999999999999999999999991) = -3.9086503371292664488601602702496216E-32
--		x"0000000000000000000000000000000039"); -- LUT(33) = log10 (0.999999999999999999999999999999991) = -3.9086503371292664488601602702494633E-33
--


-- ====== FIN declaraci�n
-- declaracion de meomria de ln para la parte de x>1

-- ====== Comienzo declaraci�n
-- declaracion de meomria de ln para la parte de x<1

type mlut_LogShN is array (0 to P-1) of std_logic_vector (4*P-1 downto 0);
-- los resultados est�n normalizados en 0.yyyyyyy (para precisi�n 7),
-- en 0.yyyyyyyyyyyyyyyy (para precisi�n 16)
-- en 0.yyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyy (para precisi�n 34)

signal lut_Log10ShN9: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"0413926", -- LUT(1) = log10 (1.1) = 0.041392685
		x"0043213", -- LUT(2) = log10 (1.01) = 0.0043213738
		x"0004340", -- LUT(3) = log10 (1.001) = 0.00043407748
		x"0000434", -- LUT(4) = log10 (1.0001) = 0.000043427277
		x"0000043", -- LUT(5) = log10 (1.00001) = 0.0000043429231
		x"0000004"); -- LUT(6) = log10 (1.000001) = 4.3429426E-7

signal lut_Log10ShN8: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"0791812", -- LUT(1) = log10 (1.2) = 0.079181246
		x"0086001", -- LUT(2) = log10 (1.02) = 0.0086001718
		x"0008677", -- LUT(3) = log10 (1.002) = 0.00086772153
		x"0000868", -- LUT(4) = log10 (1.0002) = 0.000086850212
		x"0000086", -- LUT(5) = log10 (1.00002) = 0.0000086858028
		x"0000008"); -- LUT(6) = log10 (1.000002) = 8.6858810E-7

signal lut_Log10ShN7: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"1139433", -- LUT(1) = log10 (1.3) = 0.11394335
		x"0128372", -- LUT(2) = log10 (1.03) = 0.012837225
		x"0013009", -- LUT(3) = log10 (1.003) = 0.0013009330
		x"0001302", -- LUT(4) = log10 (1.0003) = 0.00013026881
		x"0000130", -- LUT(5) = log10 (1.00003) = 0.000013028639
		x"0000013"); -- LUT(6) = log10 (1.000003) = 0.0000013028815

signal lut_Log10ShN6: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"1461280", -- LUT(1) = log10 (1.4) = 0.14612804
		x"0170333", -- LUT(2) = log10 (1.04) = 0.017033339
		x"0017337", -- LUT(3) = log10 (1.004) = 0.0017337128
		x"0001736", -- LUT(4) = log10 (1.0004) = 0.00017368306
		x"0000173", -- LUT(5) = log10 (1.00004) = 0.000017371432
		x"0000017"); -- LUT(6) = log10 (1.000004) = 0.0000017371745

signal lut_Log10ShN5: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"1760912", -- LUT(1) = log10 (1.5) = 0.17609126
		x"0211892", -- LUT(2) = log10 (1.05) = 0.021189299
		x"0021660", -- LUT(3) = log10 (1.005) = 0.0021660618
		x"0002170", -- LUT(4) = log10 (1.0005) = 0.00021709297
		x"0000217", -- LUT(5) = log10 (1.00005) = 0.000021714181
		x"0000021"); -- LUT(6) = log10 (1.000005) = 0.0000021714670

signal lut_Log10ShN4: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"2041199", -- LUT(1) = log10 (1.6) = 0.20411998
		x"0253058", -- LUT(2) = log10 (1.06) = 0.025305865
		x"0025979", -- LUT(3) = log10 (1.006) = 0.0025979807
		x"0002604", -- LUT(4) = log10 (1.0006) = 0.00026049855
		x"0000260", -- LUT(5) = log10 (1.00006) = 0.000026056887
		x"0000026"); -- LUT(6) = log10 (1.000006) = 0.0000026057591

signal lut_Log10ShN3: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"2304489", -- LUT(1) = log10 (1.7) = 0.23044892
		x"0293837", -- LUT(2) = log10 (1.07) = 0.029383778
		x"0030294", -- LUT(3) = log10 (1.007) = 0.0030294706
		x"0003038", -- LUT(4) = log10 (1.0007) = 0.00030389978
		x"0000303", -- LUT(5) = log10 (1.00007) = 0.000030399550
		x"0000030"); -- LUT(6) = log10 (1.000007) = 0.0000030400507

signal lut_Log10ShN2: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"2552725", -- LUT(1) = log10 (1.8) = 0.25527251
		x"0334237", -- LUT(2) = log10 (1.08) = 0.033423755
		x"0034605", -- LUT(3) = log10 (1.008) = 0.0034605321
		x"0003472", -- LUT(4) = log10 (1.0008) = 0.00034729669
		x"0000347", -- LUT(5) = log10 (1.00008) = 0.000034742169
		x"0000034"); -- LUT(6) = log10 (1.000008) = 0.0000034743420

signal lut_Log10ShN1: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"2787536", -- LUT(1) = log10 (1.9) = 0.27875360
		x"0374264", -- LUT(2) = log10 (1.09) = 0.037426498
		x"0038911", -- LUT(3) = log10 (1.009) = 0.0038911662
		x"0003906", -- LUT(4) = log10 (1.0009) = 0.00039068925
		x"0000390", -- LUT(5) = log10 (1.00009) = 0.000039084745
		x"0000039"); -- LUT(6) = log10 (1.000009) = 0.0000039086327

signal lut_Log10ShN0: mlut_LogShN := (
		x"0000000", -- LUT(0), No usada
		x"3010300", -- LUT(1) = log10 (2.0) = 0.30103000
		x"0413926", -- LUT(2) = log10 (1.10) = 0.041392685
		x"0043213", -- LUT(3) = log10 (1.010) = 0.0043213738
		x"0004340", -- LUT(4) = log10 (1.0010) = 0.00043407748
		x"0000434", -- LUT(5) = log10 (1.00010) = 0.000043427277
		x"0000043"); -- LUT(6) = log10 (1.000010) = 0.0000043429231
--
--
--signal lut_Log10ShN9: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"0413926851582250", -- LUT(1) = log10 (1.1) = 0.041392685158225041
--		x"0043213737826425", -- LUT(2) = log10 (1.01) = 0.0043213737826425743
--		x"0004340774793186", -- LUT(3) = log10 (1.001) = 0.00043407747931864067
--		x"0000434272768626", -- LUT(4) = log10 (1.0001) = 0.000043427276862669637
--		x"0000043429231044", -- LUT(5) = log10 (1.00001) = 0.0000043429231044531869
--		x"0000004342942647", -- LUT(6) = log10 (1.000001) = 4.3429426475615564E-7
--		x"0000000434294460", -- LUT(7) = log10 (1.0000001) = 4.3429446018852918E-8
--		x"0000000043429447", -- LUT(8) = log10 (1.00000001) = 4.3429447973177943E-9
--		x"0000000004342944", -- LUT(9) = log10 (1.000000001) = 4.3429448168610459E-10
--		x"0000000000434294", -- LUT(10) = log10 (1.0000000001) = 4.3429448188153710E-11
--		x"0000000000043429", -- LUT(11) = log10 (1.00000000001) = 4.3429448190108036E-12
--		x"0000000000004342", -- LUT(12) = log10 (1.000000000001) = 4.3429448190303468E-13
--		x"0000000000000434", -- LUT(13) = log10 (1.0000000000001) = 4.3429448190323011E-14
--		x"0000000000000043", -- LUT(14) = log10 (1.00000000000001) = 4.3429448190324966E-15
--		x"0000000000000004"); -- LUT(15) = log10 (1.000000000000001) = 4.3429448190325161E-16
--
--signal lut_Log10ShN8: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"0791812460476248", -- LUT(1) = log10 (1.2) = 0.079181246047624828
--		x"0086001717619175", -- LUT(2) = log10 (1.02) = 0.0086001717619175610
--		x"0008677215312269", -- LUT(3) = log10 (1.002) = 0.00086772153122691249
--		x"0000868502116489", -- LUT(4) = log10 (1.0002) = 0.000086850211648957229
--		x"0000086858027803", -- LUT(5) = log10 (1.00002) = 0.0000086858027803267571
--		x"0000008685880952", -- LUT(6) = log10 (1.000002) = 8.6858809521869797E-7
--		x"0000000868588876", -- LUT(7) = log10 (1.0000002) = 8.6858887694761886E-8
--		x"0000000086858895", -- LUT(8) = log10 (1.00000002) = 8.6858895512061413E-9
--		x"0000000008685889", -- LUT(9) = log10 (1.000000002) = 8.6858896293791469E-10
--		x"0000000000868588", -- LUT(10) = log10 (1.0000000002) = 8.6858896371964476E-11
--		x"0000000000086858", -- LUT(11) = log10 (1.00000000002) = 8.6858896379781777E-12
--		x"0000000000008685", -- LUT(12) = log10 (1.000000000002) = 8.6858896380563507E-13
--		x"0000000000000868", -- LUT(13) = log10 (1.0000000000002) = 8.6858896380641680E-14
--		x"0000000000000086", -- LUT(14) = log10 (1.00000000000002) = 8.6858896380649497E-15
--		x"0000000000000008"); -- LUT(15) = log10 (1.000000000000002) = 8.6858896380650279E-16
--
--signal lut_Log10ShN7: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"1139433523068367", -- LUT(1) = log10 (1.3) = 0.11394335230683677
--		x"0128372247051722", -- LUT(2) = log10 (1.03) = 0.012837224705172205
--		x"0013009330204181", -- LUT(3) = log10 (1.003) = 0.0013009330204181188
--		x"0001302688052270", -- LUT(4) = log10 (1.0003) = 0.00013026880522706100
--		x"0000130286390284", -- LUT(5) = log10 (1.00003) = 0.000013028639028489261
--		x"0000013028814913", -- LUT(6) = log10 (1.000003) = 0.0000013028814913884956
--		x"0000001302883250", -- LUT(7) = log10 (1.0000003) = 1.3028832502772777E-7
--		x"0000000130288342", -- LUT(8) = log10 (1.00000003) = 1.3028834261665042E-8
--		x"0000000013028834", -- LUT(9) = log10 (1.000000003) = 1.3028834437554303E-9
--		x"0000000001302883", -- LUT(10) = log10 (1.0000000003) = 1.3028834455143230E-10
--		x"0000000000130288", -- LUT(11) = log10 (1.00000000003) = 1.3028834456902122E-11
--		x"0000000000013028", -- LUT(12) = log10 (1.000000000003) = 1.3028834457078012E-12
--		x"0000000000001302", -- LUT(13) = log10 (1.0000000000003) = 1.3028834457095601E-13
--		x"0000000000000130", -- LUT(14) = log10 (1.00000000000003) = 1.3028834457097359E-14
--		x"0000000000000013"); -- LUT(15) = log10 (1.000000000000003) = 1.3028834457097535E-15
--
--signal lut_Log10ShN6: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"1461280356782380", -- LUT(1) = log10 (1.4) = 0.14612803567823803
--		x"0170333392987803", -- LUT(2) = log10 (1.04) = 0.017033339298780355
--		x"0017337128090005", -- LUT(3) = log10 (1.004) = 0.0017337128090005298
--		x"0001736830584649", -- LUT(4) = log10 (1.0004) = 0.00017368305846491882
--		x"0000173714318498", -- LUT(5) = log10 (1.00004) = 0.000017371431849809222
--		x"0000017371744532", -- LUT(6) = log10 (1.000004) = 0.0000017371744532664170
--		x"0000001737177580", -- LUT(7) = log10 (1.0000004) = 1.7371775801775144E-7
--		x"0000000173717789", -- LUT(8) = log10 (1.00000004) = 1.7371778928694497E-8
--		x"0000000017371779", -- LUT(9) = log10 (1.000000004) = 1.7371779241386515E-9
--		x"0000000001737177", -- LUT(10) = log10 (1.0000000004) = 1.7371779272655717E-10
--		x"0000000000173717", -- LUT(11) = log10 (1.00000000004) = 1.7371779275782638E-11
--		x"0000000000017371", -- LUT(12) = log10 (1.000000000004) = 1.7371779276095330E-12
--		x"0000000000001737", -- LUT(13) = log10 (1.0000000000004) = 1.7371779276126599E-13
--		x"0000000000000173", -- LUT(14) = log10 (1.00000000000004) = 1.7371779276129726E-14
--		x"0000000000000017"); -- LUT(15) = log10 (1.000000000000004) = 1.7371779276130038E-15
--
--signal lut_Log10ShN5: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"1760912590556812", -- LUT(1) = log10 (1.5) = 0.17609125905568124
--		x"0211892990699380", -- LUT(2) = log10 (1.05) = 0.021189299069938073
--		x"0021660617565076", -- LUT(3) = log10 (1.005) = 0.0021660617565076762
--		x"0002170929722302", -- LUT(4) = log10 (1.0005) = 0.00021709297223020828
--		x"0000217141812451", -- LUT(5) = log10 (1.00005) = 0.000021714181245155137
--		x"0000021714669808", -- LUT(6) = log10 (1.000005) = 0.0000021714669808533309
--		x"0000002171471866", -- LUT(7) = log10 (1.0000005) = 2.1714718666483377E-7
--		x"0000000217147235", -- LUT(8) = log10 (1.00000005) = 2.1714723552294507E-8
--		x"0000000021714724", -- LUT(9) = log10 (1.000000005) = 2.1714724040875781E-9
--		x"0000000002171472", -- LUT(10) = log10 (1.0000000005) = 2.1714724089733910E-10
--		x"0000000000217147", -- LUT(11) = log10 (1.00000000005) = 2.1714724094619723E-11
--		x"0000000000021714", -- LUT(12) = log10 (1.000000000005) = 2.1714724095108305E-12
--		x"0000000000002171", -- LUT(13) = log10 (1.0000000000005) = 2.1714724095157163E-13
--		x"0000000000000217", -- LUT(14) = log10 (1.00000000000005) = 2.1714724095162049E-14
--		x"0000000000000021"); -- LUT(15) = log10 (1.000000000000005) = 2.1714724095162537E-15
--
--signal lut_Log10ShN4: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"2041199826559247", -- LUT(1) = log10 (1.6) = 0.20411998265592478
--		x"0253058652647702", -- LUT(2) = log10 (1.06) = 0.025305865264770241
--		x"0025979807199085", -- LUT(3) = log10 (1.006) = 0.0025979807199085923
--		x"0002604985473903", -- LUT(4) = log10 (1.0006) = 0.00026049854739034682
--		x"0000260568872153", -- LUT(5) = log10 (1.00006) = 0.000026056887215395479
--		x"0000026057590741", -- LUT(6) = log10 (1.000006) = 0.0000026057590741501058
--		x"0000002605766109", -- LUT(7) = log10 (1.0000006) = 2.6057661096897562E-7
--		x"0000000260576681", -- LUT(8) = log10 (1.00000006) = 2.6057668132465074E-8
--		x"0000000026057668", -- LUT(9) = log10 (1.000000006) = 2.6057668836022103E-9
--		x"0000000002605766", -- LUT(10) = log10 (1.0000000006) = 2.6057668906377809E-10
--		x"0000000000260576", -- LUT(11) = log10 (1.00000000006) = 2.6057668913413380E-11
--		x"0000000000026057", -- LUT(12) = log10 (1.000000000006) = 2.6057668914116937E-12
--		x"0000000000002605", -- LUT(13) = log10 (1.0000000000006) = 2.6057668914187292E-13
--		x"0000000000000260", -- LUT(14) = log10 (1.00000000000006) = 2.6057668914194328E-14
--		x"0000000000000026"); -- LUT(15) = log10 (1.000000000000006) = 2.6057668914195031E-15
--
--signal lut_Log10ShN3: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"2304489213782739", -- LUT(1) = log10 (1.7) = 0.23044892137827393
--		x"0293837776852096", -- LUT(2) = log10 (1.07) = 0.029383777685209641
--		x"0030294705536180", -- LUT(3) = log10 (1.007) = 0.0030294705536180072
--		x"0003038997848124", -- LUT(4) = log10 (1.0007) = 0.00030389978481249181
--		x"0000303995497613", -- LUT(5) = log10 (1.00007) = 0.000030399549761398694
--		x"0000030400507331", -- LUT(6) = log10 (1.000007) = 0.0000030400507331576102
--		x"0000003040060309", -- LUT(7) = log10 (1.0000007) = 3.0400603093017787E-7
--		x"0000000304006126", -- LUT(8) = log10 (1.00000007) = 3.0400612669206197E-8
--		x"0000000030400613", -- LUT(9) = log10 (1.000000007) = 3.0400613626825480E-9
--		x"0000000003040061", -- LUT(10) = log10 (1.0000000007) = 3.0400613722587413E-10
--		x"0000000000304006", -- LUT(11) = log10 (1.00000000007) = 3.0400613732163606E-11
--		x"0000000000030400", -- LUT(12) = log10 (1.000000000007) = 3.0400613733121226E-12
--		x"0000000000003040", -- LUT(13) = log10 (1.0000000000007) = 3.0400613733216988E-13
--		x"0000000000000304", -- LUT(14) = log10 (1.00000000000007) = 3.0400613733226564E-14
--		x"0000000000000030"); -- LUT(15) = log10 (1.000000000000007) = 3.0400613733227522E-15
--
--signal lut_Log10ShN2: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"2552725051033060", -- LUT(1) = log10 (1.8) = 0.25527250510330607
--		x"0334237554869497", -- LUT(2) = log10 (1.08) = 0.033423755486949702
--		x"0034605321095064", -- LUT(3) = log10 (1.008) = 0.0034605321095064862
--		x"0003472966853635", -- LUT(4) = log10 (1.0008) = 0.00034729668536354069
--		x"0000347421688840", -- LUT(5) = log10 (1.00008) = 0.000034742168884033200
--		x"0000034743419578", -- LUT(6) = log10 (1.000008) = 0.0000034743419578767129
--		x"0000003474354465", -- LUT(7) = log10 (1.0000008) = 3.4743544654844137E-7
--		x"0000000347435571", -- LUT(8) = log10 (1.00000008) = 3.4743557162517878E-8
--		x"0000000034743558", -- LUT(9) = log10 (1.000000008) = 3.4743558413285913E-9
--		x"0000000003474355", -- LUT(10) = log10 (1.0000000008) = 3.4743558538362723E-10
--		x"0000000000347435", -- LUT(11) = log10 (1.00000000008) = 3.4743558550870404E-11
--		x"0000000000034743", -- LUT(12) = log10 (1.000000000008) = 3.4743558552121172E-12
--		x"0000000000003474", -- LUT(13) = log10 (1.0000000000008) = 3.4743558552246249E-13
--		x"0000000000000347", -- LUT(14) = log10 (1.00000000000008) = 3.4743558552258756E-14
--		x"0000000000000034"); -- LUT(15) = log10 (1.000000000000008) = 3.4743558552260007E-15
--
--signal lut_Log10ShN1: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"2787536009528289", -- LUT(1) = log10 (1.9) = 0.27875360095282896
--		x"0374264979406236", -- LUT(2) = log10 (1.09) = 0.037426497940623635
--		x"0038911662369105", -- LUT(3) = log10 (1.009) = 0.0038911662369105217
--		x"0003906892499101", -- LUT(4) = log10 (1.0009) = 0.00039068924991013103
--		x"0000390847445841", -- LUT(5) = log10 (1.00009) = 0.000039084744584167392
--		x"0000039086327483", -- LUT(6) = log10 (1.000009) = 0.0000039086327483082822
--		x"0000003908648578", -- LUT(7) = log10 (1.0000009) = 3.9086485782376701E-7
--		x"0000000390865016", -- LUT(8) = log10 (1.00000009) = 3.9086501612400118E-8
--		x"0000000039086503", -- LUT(9) = log10 (1.000000009) = 3.9086503195403400E-9
--		x"0000000003908650", -- LUT(10) = log10 (1.0000000009) = 3.9086503353703738E-10
--		x"0000000000390865", -- LUT(11) = log10 (1.00000000009) = 3.9086503369533772E-11
--		x"0000000000039086", -- LUT(12) = log10 (1.000000000009) = 3.9086503371116775E-12
--		x"0000000000003908", -- LUT(13) = log10 (1.0000000000009) = 3.9086503371275076E-13
--		x"0000000000000390", -- LUT(14) = log10 (1.00000000000009) = 3.9086503371290906E-14
--		x"0000000000000039"); -- LUT(15) = log10 (1.000000000000009) = 3.9086503371292489E-15
--
--signal lut_Log10ShN0: mlut_LogShN := (
--		x"0000000000000000", -- LUT(0), No usada
--		x"3010299956639812", -- LUT(1) = log10 (2.0) = 0.30102999566398120
--		x"0413926851582250", -- LUT(2) = log10 (1.10) = 0.041392685158225041
--		x"0043213737826425", -- LUT(3) = log10 (1.010) = 0.0043213737826425743
--		x"0004340774793186", -- LUT(4) = log10 (1.0010) = 0.00043407747931864067
--		x"0000434272768626", -- LUT(5) = log10 (1.00010) = 0.000043427276862669637
--		x"0000043429231044", -- LUT(6) = log10 (1.000010) = 0.0000043429231044531869
--		x"0000004342942647", -- LUT(7) = log10 (1.0000010) = 4.3429426475615564E-7
--		x"0000000434294460", -- LUT(8) = log10 (1.00000010) = 4.3429446018852918E-8
--		x"0000000043429447", -- LUT(9) = log10 (1.000000010) = 4.3429447973177943E-9
--		x"0000000004342944", -- LUT(10) = log10 (1.0000000010) = 4.3429448168610459E-10
--		x"0000000000434294", -- LUT(11) = log10 (1.00000000010) = 4.3429448188153710E-11
--		x"0000000000043429", -- LUT(12) = log10 (1.000000000010) = 4.3429448190108036E-12
--		x"0000000000004342", -- LUT(13) = log10 (1.0000000000010) = 4.3429448190303468E-13
--		x"0000000000000434", -- LUT(14) = log10 (1.00000000000010) = 4.3429448190323011E-14
--		x"0000000000000043"); -- LUT(15) = log10 (1.000000000000010) = 4.3429448190324966E-15
--
--signal lut_Log10ShN9: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"0413926851582250407501999712430242", -- LUT(1) = log10 (1.1) = 0.041392685158225040750199971243024242
--		x"0043213737826425742751881782229379", -- LUT(2) = log10 (1.01) = 0.0043213737826425742751881782229379132
--		x"0004340774793186406689213877779888", -- LUT(3) = log10 (1.001) = 0.00043407747931864066892138777798886602
--		x"0000434272768626696373135275850982", -- LUT(4) = log10 (1.0001) = 0.000043427276862669637313527585098268131
--		x"0000043429231044531868554934716343", -- LUT(5) = log10 (1.00001) = 0.0000043429231044531868554934716343971840
--		x"0000004342942647561556407439426436", -- LUT(6) = log10 (1.000001) = 4.3429426475615564074394264367770704E-7
--		x"0000000434294460188529180136701973", -- LUT(7) = log10 (1.0000001) = 4.3429446018852918013670197358779472E-8
--		x"0000000043429447973177943261135240", -- LUT(8) = log10 (1.00000001) = 4.3429447973177943261135240219573514E-9
--		x"0000000004342944816861045868442678", -- LUT(9) = log10 (1.000000001) = 4.3429448168610458684426783228355094E-10
--		x"0000000000434294481881537103557413", -- LUT(10) = log10 (1.0000000001) = 4.3429448188153710355741397580695090E-11
--		x"0000000000043429448190108035524162", -- LUT(11) = log10 (1.00000000001) = 4.3429448190108035524162713626107944E-12
--		x"0000000000004342944819030346804101", -- LUT(12) = log10 (1.000000000001) = 4.3429448190303468041017743776760682E-13
--		x"0000000000000434294481903230112927", -- LUT(13) = log10 (1.0000000000001) = 4.3429448190323011292703375777287080E-14
--		x"0000000000000043429448190324965617", -- LUT(14) = log10 (1.00000000000001) = 4.3429448190324965617871940267194331E-15
--		x"0000000000000004342944819032516105", -- LUT(15) = log10 (1.000000000000001) = 4.3429448190325161050388796729083602E-16
--		x"0000000000000000434294481903251805", -- LUT(16) = log10 (1.0000000000000001) = 4.3429448190325180593640482375401515E-17
--		x"0000000000000000043429448190325182", -- LUT(17) = log10 (1.00000000000000001) = 4.3429448190325182547965650940034596E-18
--		x"0000000000000000004342944819032518", -- LUT(18) = log10 (1.000000000000000001) = 4.3429448190325182743398167796497917E-19
--		x"0000000000000000000434294481903251", -- LUT(19) = log10 (1.0000000000000000001) = 4.3429448190325182762941419482144249E-20
--		x"0000000000000000000043429448190325", -- LUT(20) = log10 (1.00000000000000000001) = 4.3429448190325182764895744650708882E-21
--		x"0000000000000000000004342944819032", -- LUT(21) = log10 (1.000000000000000000001) = 4.3429448190325182765091177167565346E-22
--		x"0000000000000000000000434294481903", -- LUT(22) = log10 (1.0000000000000000000001) = 4.3429448190325182765110720419250992E-23
--		x"0000000000000000000000043429448190", -- LUT(23) = log10 (1.00000000000000000000001) = 4.3429448190325182765112674744419557E-24
--		x"0000000000000000000000004342944819", -- LUT(24) = log10 (1.000000000000000000000001) = 4.3429448190325182765112870176936413E-25
--		x"0000000000000000000000000434294481", -- LUT(25) = log10 (1.0000000000000000000000001) = 4.3429448190325182765112889720188099E-26
--		x"0000000000000000000000000043429448", -- LUT(26) = log10 (1.00000000000000000000000001) = 4.3429448190325182765112891674513267E-27
--		x"0000000000000000000000000004342944", -- LUT(27) = log10 (1.000000000000000000000000001) = 4.3429448190325182765112891869945784E-28
--		x"0000000000000000000000000000434294", -- LUT(28) = log10 (1.0000000000000000000000000001) = 4.3429448190325182765112891889489036E-29
--		x"0000000000000000000000000000043429", -- LUT(29) = log10 (1.00000000000000000000000000001) = 4.3429448190325182765112891891443361E-30
--		x"0000000000000000000000000000004342", -- LUT(30) = log10 (1.000000000000000000000000000001) = 4.3429448190325182765112891891638794E-31
--		x"0000000000000000000000000000000434", -- LUT(31) = log10 (1.0000000000000000000000000000001) = 4.3429448190325182765112891891658337E-32
--		x"0000000000000000000000000000000043", -- LUT(32) = log10 (1.00000000000000000000000000000001) = 4.3429448190325182765112891891660291E-33
--		x"0000000000000000000000000000000004"); -- LUT(33) = log10 (1.000000000000000000000000000000001) = 4.3429448190325182765112891891660487E-34
--
--signal lut_Log10ShN8: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"0791812460476248277225056927041013", -- LUT(1) = log10 (1.2) = 0.079181246047624827722505692704101363
--		x"0086001717619175610489366923079453", -- LUT(2) = log10 (1.02) = 0.0086001717619175610489366923079453660
--		x"0008677215312269124928427079000758", -- LUT(3) = log10 (1.002) = 0.00086772153122691249284270790007587043
--		x"0000868502116489572288997981622109", -- LUT(4) = log10 (1.0002) = 0.000086850211648957228899798162210906629
--		x"0000086858027803267571495643873989", -- LUT(5) = log10 (1.00002) = 0.0000086858027803267571495643873989012427
--		x"0000008685880952186979656798360589", -- LUT(6) = log10 (1.000002) = 8.6858809521869796567983605898281975E-7
--		x"0000000868588876947618855836339216", -- LUT(7) = log10 (1.0000002) = 8.6858887694761885583633921667316583E-8
--		x"0000000086858895512061413304908138", -- LUT(8) = log10 (1.00000002) = 8.6858895512061413304908138849988601E-9
--		x"0000000008685889629379146926538727", -- LUT(9) = log10 (1.000000002) = 8.6858896293791469265387279920244594E-10
--		x"0000000000868588963719644758933188", -- LUT(10) = log10 (1.0000000002) = 8.6858896371964475893318865848533392E-11
--		x"0000000000086858896379781776566430", -- LUT(11) = log10 (1.00000000002) = 8.6858896379781776566430861314202672E-12
--		x"0000000000008685889638056350663384", -- LUT(12) = log10 (1.000000000002) = 8.6858896380563506633845249229652631E-13
--		x"0000000000000868588963806416796405", -- LUT(13) = log10 (1.0000000000002) = 8.6858896380641679640587719904886612E-14
--		x"0000000000000086858896380649496941", -- LUT(14) = log10 (1.00000000000002) = 8.6858896380649496941261977291246900E-15
--		x"0000000000000008685889638065027867", -- LUT(15) = log10 (1.000000000000002) = 8.6858896380650278671329403133071298E-16
--		x"0000000000000000868588963806503568", -- LUT(16) = log10 (1.0000000000000002) = 8.6858896380650356844336145718285622E-17
--		x"0000000000000000086858896380650364", -- LUT(17) = log10 (1.00000000000000002) = 8.6858896380650364661636819976817373E-18
--		x"0000000000000000008685889638065036", -- LUT(18) = log10 (1.000000000000000002) = 8.6858896380650365443366887402670651E-19
--		x"0000000000000000000868588963806503", -- LUT(19) = log10 (1.0000000000000000002) = 8.6858896380650365521539894145255980E-20
--		x"0000000000000000000086858896380650", -- LUT(20) = log10 (1.00000000000000000002) = 8.6858896380650365529357194819514513E-21
--		x"0000000000000000000008685889638065", -- LUT(21) = log10 (1.000000000000000000002) = 8.6858896380650365530138924886940366E-22
--		x"0000000000000000000000868588963806", -- LUT(22) = log10 (1.0000000000000000000002) = 8.6858896380650365530217097893682951E-23
--		x"0000000000000000000000086858896380", -- LUT(23) = log10 (1.00000000000000000000002) = 8.6858896380650365530224915194357210E-24
--		x"0000000000000000000000008685889638", -- LUT(24) = log10 (1.000000000000000000000002) = 8.6858896380650365530225696924424636E-25
--		x"0000000000000000000000000868588963", -- LUT(25) = log10 (1.0000000000000000000000002) = 8.6858896380650365530225775097431378E-26
--		x"0000000000000000000000000086858896", -- LUT(26) = log10 (1.00000000000000000000000002) = 8.6858896380650365530225782914732053E-27
--		x"0000000000000000000000000008685889", -- LUT(27) = log10 (1.000000000000000000000000002) = 8.6858896380650365530225783696462120E-28
--		x"0000000000000000000000000000868588", -- LUT(28) = log10 (1.0000000000000000000000000002) = 8.6858896380650365530225783774635127E-29
--		x"0000000000000000000000000000086858", -- LUT(29) = log10 (1.00000000000000000000000000002) = 8.6858896380650365530225783782452427E-30
--		x"0000000000000000000000000000008685", -- LUT(30) = log10 (1.000000000000000000000000000002) = 8.6858896380650365530225783783234158E-31
--		x"0000000000000000000000000000000868", -- LUT(31) = log10 (1.0000000000000000000000000000002) = 8.6858896380650365530225783783312331E-32
--		x"0000000000000000000000000000000086", -- LUT(32) = log10 (1.00000000000000000000000000000002) = 8.6858896380650365530225783783320148E-33
--		x"0000000000000000000000000000000008"); -- LUT(33) = log10 (1.000000000000000000000000000000002) = 8.6858896380650365530225783783320930E-34
--
--signal lut_Log10ShN7: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"1139433523068367692065051579423284", -- LUT(1) = log10 (1.3) = 0.11394335230683676920650515794232843
--		x"0128372247051722051710711945802394", -- LUT(2) = log10 (1.03) = 0.012837224705172205171071194580239424
--		x"0013009330204181188008262788634812", -- LUT(3) = log10 (1.003) = 0.0013009330204181188008262788634812689
--		x"0001302688052270610037808717292515", -- LUT(4) = log10 (1.0003) = 0.00013026880522706100378087172925158811
--		x"0000130286390284892607608187240164", -- LUT(5) = log10 (1.00003) = 0.000013028639028489260760818724016476778
--		x"0000013028814913884955598628494412", -- LUT(6) = log10 (1.000003) = 0.0000013028814913884955598628494412367446
--		x"0000001302883250277277712984641145", -- LUT(7) = log10 (1.0000003) = 1.3028832502772777129846411452584201E-7
--		x"0000000130288342616650418817207943", -- LUT(8) = log10 (1.00000003) = 1.3028834261665041881720794309126113E-8
--		x"0000000013028834437554303182974038", -- LUT(9) = log10 (1.000000003) = 1.3028834437554303182974038606545383E-9
--		x"0000000001302883445514322966136009", -- LUT(10) = log10 (1.0000000003) = 1.3028834455143229661360099376693054E-10
--		x"0000000000130288344569021223126813", -- LUT(11) = log10 (1.00000000003) = 1.3028834456902122312681312895392186E-11
--		x"0000000000013028834457078011577848", -- LUT(12) = log10 (1.000000000003) = 1.3028834457078011577848260321757223E-12
--		x"0000000000001302883445709560050436", -- LUT(13) = log10 (1.0000000000003) = 1.3028834457095600504365303325138756E-13
--		x"0000000000000130288344570973593970", -- LUT(14) = log10 (1.00000000000003) = 1.3028834457097359397017011108084360E-14
--		x"0000000000000013028834457097535286", -- LUT(15) = log10 (1.000000000000003) = 1.3028834457097535286282181921204995E-15
--		x"0000000000000001302883445709755287", -- LUT(16) = log10 (1.0000000000000003) = 1.3028834457097552875208699002865319E-16
--		x"0000000000000000130288344570975546", -- LUT(17) = log10 (1.00000000000000003) = 1.3028834457097554634101350711034834E-17
--		x"0000000000000000013028834457097554", -- LUT(18) = log10 (1.000000000000000003) = 1.3028834457097554809990615881851820E-18
--		x"0000000000000000001302883445709755", -- LUT(19) = log10 (1.0000000000000000003) = 1.3028834457097554827579542398933519E-19
--		x"0000000000000000000130288344570975", -- LUT(20) = log10 (1.00000000000000000003) = 1.3028834457097554829338435050641689E-20
--		x"0000000000000000000013028834457097", -- LUT(21) = log10 (1.000000000000000000003) = 1.3028834457097554829514324315812506E-21
--		x"0000000000000000000001302883445709", -- LUT(22) = log10 (1.0000000000000000000003) = 1.3028834457097554829531913242329588E-22
--		x"0000000000000000000000130288344570", -- LUT(23) = log10 (1.00000000000000000000003) = 1.3028834457097554829533672134981296E-23
--		x"0000000000000000000000013028834457", -- LUT(24) = log10 (1.000000000000000000000003) = 1.3028834457097554829533848024246467E-24
--		x"0000000000000000000000001302883445", -- LUT(25) = log10 (1.0000000000000000000000003) = 1.3028834457097554829533865613172984E-25
--		x"0000000000000000000000000130288344", -- LUT(26) = log10 (1.00000000000000000000000003) = 1.3028834457097554829533867372065636E-26
--		x"0000000000000000000000000013028834", -- LUT(27) = log10 (1.000000000000000000000000003) = 1.3028834457097554829533867547954901E-27
--		x"0000000000000000000000000001302883", -- LUT(28) = log10 (1.0000000000000000000000000003) = 1.3028834457097554829533867565543827E-28
--		x"0000000000000000000000000000130288", -- LUT(29) = log10 (1.00000000000000000000000000003) = 1.3028834457097554829533867567302720E-29
--		x"0000000000000000000000000000013028", -- LUT(30) = log10 (1.000000000000000000000000000003) = 1.3028834457097554829533867567478609E-30
--		x"0000000000000000000000000000001302", -- LUT(31) = log10 (1.0000000000000000000000000000003) = 1.3028834457097554829533867567496198E-31
--		x"0000000000000000000000000000000130", -- LUT(32) = log10 (1.00000000000000000000000000000003) = 1.3028834457097554829533867567497957E-32
--		x"0000000000000000000000000000000013"); -- LUT(33) = log10 (1.000000000000000000000000000000003) = 1.3028834457097554829533867567498133E-33
--
--signal lut_Log10ShN6: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"1461280356782380259259551533171292", -- LUT(1) = log10 (1.4) = 0.14612803567823802592595515331712922
--		x"0170333392987803548477218421158075", -- LUT(2) = log10 (1.04) = 0.017033339298780354847721842115807511
--		x"0017337128090005297680271061558901", -- LUT(3) = log10 (1.004) = 0.0017337128090005297680271061558901354
--		x"0001736830584649188226381531744882", -- LUT(4) = log10 (1.0004) = 0.00017368305846491882263815317448820233
--		x"0000173714318498092215122780446167", -- LUT(5) = log10 (1.00004) = 0.000017371431849809221512278044616760358
--		x"0000017371744532664170057424059403", -- LUT(6) = log10 (1.000004) = 0.0000017371744532664170057424059403635925
--		x"0000001737177580177514437464731410", -- LUT(7) = log10 (1.0000004) = 1.7371775801775144374647314105390573E-7
--		x"0000000173717789286944968483923639", -- LUT(8) = log10 (1.00000004) = 1.7371778928694496848392363956673868E-8
--		x"0000000017371779241386514646434499", -- LUT(9) = log10 (1.000000004) = 1.7371779241386514646434499739319145E-9
--		x"0000000001737177927265571725174563", -- LUT(10) = log10 (1.0000000004) = 1.7371779272655717251745637029904161E-10
--		x"0000000000173717792757826375205318", -- LUT(11) = log10 (1.00000000004) = 1.7371779275782637520531820243490292E-11
--		x"0000000000017371779276095329547492", -- LUT(12) = log10 (1.000000000004) = 1.7371779276095329547492989259941585E-12
--		x"0000000000001737177927612659875018", -- LUT(13) = log10 (1.0000000000004) = 1.7371779276126598750189931668537889E-13
--		x"0000000000000173717792761297256704", -- LUT(14) = log10 (1.00000000000004) = 1.7371779276129725670459634164467031E-14
--		x"0000000000000017371779276130038362", -- LUT(15) = log10 (1.000000000000004) = 1.7371779276130038362486604496610641E-15
--		x"0000000000000001737177927613006963", -- LUT(16) = log10 (1.0000000000000004) = 1.7371779276130069631689301530650509E-16
--		x"0000000000000000173717792761300727", -- LUT(17) = log10 (1.00000000000000004) = 1.7371779276130072758609571234062750E-17
--		x"0000000000000000017371779276130073", -- LUT(18) = log10 (1.000000000000000004) = 1.7371779276130073071301598204404057E-18
--		x"0000000000000000001737177927613007", -- LUT(19) = log10 (1.0000000000000000004) = 1.7371779276130073102570800901438189E-19
--		x"0000000000000000000173717792761300", -- LUT(20) = log10 (1.00000000000000000004) = 1.7371779276130073105697721171141602E-20
--		x"0000000000000000000017371779276130", -- LUT(21) = log10 (1.000000000000000000004) = 1.7371779276130073106010413198111943E-21
--		x"0000000000000000000001737177927613", -- LUT(22) = log10 (1.0000000000000000000004) = 1.7371779276130073106041682400808977E-22
--		x"0000000000000000000000173717792761", -- LUT(23) = log10 (1.00000000000000000000004) = 1.7371779276130073106044809321078681E-23
--		x"0000000000000000000000017371779276", -- LUT(24) = log10 (1.000000000000000000000004) = 1.7371779276130073106045122013105651E-24
--		x"0000000000000000000000001737177927", -- LUT(25) = log10 (1.0000000000000000000000004) = 1.7371779276130073106045153282308348E-25
--		x"0000000000000000000000000173717792", -- LUT(26) = log10 (1.00000000000000000000000004) = 1.7371779276130073106045156409228618E-26
--		x"0000000000000000000000000017371779", -- LUT(27) = log10 (1.000000000000000000000000004) = 1.7371779276130073106045156721920645E-27
--		x"0000000000000000000000000001737177", -- LUT(28) = log10 (1.0000000000000000000000000004) = 1.7371779276130073106045156753189847E-28
--		x"0000000000000000000000000000173717", -- LUT(29) = log10 (1.00000000000000000000000000004) = 1.7371779276130073106045156756316768E-29
--		x"0000000000000000000000000000017371", -- LUT(30) = log10 (1.000000000000000000000000000004) = 1.7371779276130073106045156756629460E-30
--		x"0000000000000000000000000000001737", -- LUT(31) = log10 (1.0000000000000000000000000000004) = 1.7371779276130073106045156756660729E-31
--		x"0000000000000000000000000000000173", -- LUT(32) = log10 (1.00000000000000000000000000000004) = 1.7371779276130073106045156756663856E-32
--		x"0000000000000000000000000000000017"); -- LUT(33) = log10 (1.000000000000000000000000000000004) = 1.7371779276130073106045156756664169E-33
--
--signal lut_Log10ShN5: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"1760912590556812420812890085306222", -- LUT(1) = log10 (1.5) = 0.17609125905568124208128900853062228
--		x"0211892990699380727935052671232584", -- LUT(2) = log10 (1.05) = 0.021189299069938072793505267123258476
--		x"0021660617565076762304206377566908", -- LUT(3) = log10 (1.005) = 0.0021660617565076762304206377566908634
--		x"0002170929722302082819128837510668", -- LUT(4) = log10 (1.0005) = 0.00021709297223020828191288375106682338
--		x"0000217141812451551371724216752147", -- LUT(5) = log10 (1.00005) = 0.000021714181245155137172421675214706137
--		x"0000021714669808533308831621930838", -- LUT(6) = log10 (1.000005) = 0.0000021714669808533308831621930838274571
--		x"0000002171471866648337715157127899", -- LUT(7) = log10 (1.0000005) = 2.1714718666483377151571278999460754E-7
--		x"0000000217147235522945070990943954", -- LUT(8) = log10 (1.00000005) = 2.1714723552294507099094395432311094E-8
--		x"0000000021714724040875781325606000", -- LUT(9) = log10 (1.000000005) = 2.1714724040875781325606000937208942E-9
--		x"0000000002171472408973391036057535", -- LUT(10) = log10 (1.0000000005) = 2.1714724089733910360575358440776107E-10
--		x"0000000000217147240946197232801954", -- LUT(11) = log10 (1.00000000005) = 2.1714724094619723280195476764678300E-11
--		x"0000000000021714724095108304572318", -- LUT(12) = log10 (1.000000000005) = 2.1714724095108304572318720423407989E-12
--		x"0000000000002171472409515716270153", -- LUT(13) = log10 (1.0000000000005) = 2.1714724095157162701532657107544956E-13
--		x"0000000000000217147240951620485144", -- LUT(14) = log10 (1.00000000000005) = 2.1714724095162048514454066899141294E-14
--		x"0000000000000021714724095162537095", -- LUT(15) = log10 (1.000000000000005) = 2.1714724095162537095746208039532754E-15
--		x"0000000000000002171472409516258595", -- LUT(16) = log10 (1.0000000000000005) = 2.1714724095162585953875422155184218E-16
--		x"0000000000000000217147240951625908", -- LUT(17) = log10 (1.00000000000000005) = 2.1714724095162590839688343566765488E-17
--		x"0000000000000000021714724095162591", -- LUT(18) = log10 (1.000000000000000005) = 2.1714724095162591328269635707923776E-18
--		x"0000000000000000002171472409516259", -- LUT(19) = log10 (1.0000000000000000005) = 2.1714724095162591377127764922039606E-19
--		x"0000000000000000000217147240951625", -- LUT(20) = log10 (1.00000000000000000005) = 2.1714724095162591382013577843451189E-20
--		x"0000000000000000000021714724095162", -- LUT(21) = log10 (1.000000000000000000005) = 2.1714724095162591382502159135592348E-21
--		x"0000000000000000000002171472409516", -- LUT(22) = log10 (1.0000000000000000000005) = 2.1714724095162591382551017264806463E-22
--		x"0000000000000000000000217147240951", -- LUT(23) = log10 (1.00000000000000000000005) = 2.1714724095162591382555903077727875E-23
--		x"0000000000000000000000021714724095", -- LUT(24) = log10 (1.000000000000000000000005) = 2.1714724095162591382556391659020016E-24
--		x"0000000000000000000000002171472409", -- LUT(25) = log10 (1.0000000000000000000000005) = 2.1714724095162591382556440517149230E-25
--		x"0000000000000000000000000217147240", -- LUT(26) = log10 (1.00000000000000000000000005) = 2.1714724095162591382556445402962152E-26
--		x"0000000000000000000000000021714724", -- LUT(27) = log10 (1.000000000000000000000000005) = 2.1714724095162591382556445891543444E-27
--		x"0000000000000000000000000002171472", -- LUT(28) = log10 (1.0000000000000000000000000005) = 2.1714724095162591382556445940401573E-28
--		x"0000000000000000000000000000217147", -- LUT(29) = log10 (1.00000000000000000000000000005) = 2.1714724095162591382556445945287386E-29
--		x"0000000000000000000000000000021714", -- LUT(30) = log10 (1.000000000000000000000000000005) = 2.1714724095162591382556445945775967E-30
--		x"0000000000000000000000000000002171", -- LUT(31) = log10 (1.0000000000000000000000000000005) = 2.1714724095162591382556445945824825E-31
--		x"0000000000000000000000000000000217", -- LUT(32) = log10 (1.00000000000000000000000000000005) = 2.1714724095162591382556445945829711E-32
--		x"0000000000000000000000000000000021"); -- LUT(33) = log10 (1.000000000000000000000000000000005) = 2.1714724095162591382556445945830200E-33
--
--signal lut_Log10ShN4: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"2041199826559247808549555788979721", -- LUT(1) = log10 (1.6) = 0.20411998265592478085495557889797211
--		x"0253058652647702408467311863517496", -- LUT(2) = log10 (1.06) = 0.025305865264770240846731186351749619
--		x"0025979807199085923119629850040210", -- LUT(3) = log10 (1.006) = 0.0025979807199085923119629850040210818
--		x"0002604985473903468178546109174371", -- LUT(4) = log10 (1.0006) = 0.00026049854739034681785461091743713901
--		x"0000260568872153954794562288290832", -- LUT(5) = log10 (1.00006) = 0.000026056887215395479456228829083273360
--		x"0000026057590741501057693601731995", -- LUT(6) = log10 (1.000006) = 0.0000026057590741501057693601731995175785
--		x"0000002605766109689756231939742738", -- LUT(7) = log10 (1.0000006) = 2.6057661096897562319397427381882757E-7
--		x"0000000260576681324650735024157352", -- LUT(8) = log10 (1.00000006) = 2.6057668132465073502415735283042017E-8
--		x"0000000026057668836022103229174431", -- LUT(9) = log10 (1.000000006) = 2.6057668836022103229174431721020301E-9
--		x"0000000002605766890637780898793612", -- LUT(10) = log10 (1.0000000006) = 2.6057668906377808987936122505572283E-10
--		x"0000000000260576689134133795916731", -- LUT(11) = log10 (1.00000000006) = 2.6057668913413379591673151047919900E-11
--		x"0000000000026057668914116936652325", -- LUT(12) = log10 (1.000000000006) = 2.6057668914116936652325462498046071E-12
--		x"0000000000002605766891418729235839", -- LUT(13) = log10 (1.0000000000006) = 2.6057668914187292358393479729018854E-13
--		x"0000000000000260576689141943279290", -- LUT(14) = log10 (1.00000000000006) = 2.6057668914194327929000309312975736E-14
--		x"0000000000000026057668914195031486", -- LUT(15) = log10 (1.000000000000006) = 2.6057668914195031486060992549980020E-15
--		x"0000000000000002605766891419510184", -- LUT(16) = log10 (1.0000000000000006) = 2.6057668914195101841767060876466534E-16
--		x"0000000000000000260576689141951088", -- LUT(17) = log10 (1.00000000000000006) = 2.6057668914195108877337667709143046E-17
--		x"0000000000000000026057668914195109", -- LUT(18) = log10 (1.000000000000000006) = 2.6057668914195109580894728392410976E-18
--		x"0000000000000000002605766891419510", -- LUT(19) = log10 (1.0000000000000000006) = 2.6057668914195109651250434460737772E-19
--		x"0000000000000000000260576689141951", -- LUT(20) = log10 (1.00000000000000000006) = 2.6057668914195109658286005067570452E-20
--		x"0000000000000000000026057668914195", -- LUT(21) = log10 (1.000000000000000000006) = 2.6057668914195109658989562128253720E-21
--		x"0000000000000000000002605766891419", -- LUT(22) = log10 (1.0000000000000000000006) = 2.6057668914195109659059917834322046E-22
--		x"0000000000000000000000260576689141", -- LUT(23) = log10 (1.00000000000000000000006) = 2.6057668914195109659066953404928879E-23
--		x"0000000000000000000000026057668914", -- LUT(24) = log10 (1.000000000000000000000006) = 2.6057668914195109659067656961989562E-24
--		x"0000000000000000000000002605766891", -- LUT(25) = log10 (1.0000000000000000000000006) = 2.6057668914195109659067727317695631E-25
--		x"0000000000000000000000000260576689", -- LUT(26) = log10 (1.00000000000000000000000006) = 2.6057668914195109659067734353266238E-26
--		x"0000000000000000000000000026057668", -- LUT(27) = log10 (1.000000000000000000000000006) = 2.6057668914195109659067735056823298E-27
--		x"0000000000000000000000000002605766", -- LUT(28) = log10 (1.0000000000000000000000000006) = 2.6057668914195109659067735127179004E-28
--		x"0000000000000000000000000000260576", -- LUT(29) = log10 (1.00000000000000000000000000006) = 2.6057668914195109659067735134214575E-29
--		x"0000000000000000000000000000026057", -- LUT(30) = log10 (1.000000000000000000000000000006) = 2.6057668914195109659067735134918132E-30
--		x"0000000000000000000000000000002605", -- LUT(31) = log10 (1.0000000000000000000000000000006) = 2.6057668914195109659067735134988488E-31
--		x"0000000000000000000000000000000260", -- LUT(32) = log10 (1.00000000000000000000000000000006) = 2.6057668914195109659067735134995523E-32
--		x"0000000000000000000000000000000026"); -- LUT(33) = log10 (1.000000000000000000000000000000006) = 2.6057668914195109659067735134996227E-33
--
--signal lut_Log10ShN3: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"2304489213782739285401698943283370", -- LUT(1) = log10 (1.7) = 0.23044892137827392854016989432833703
--		x"0293837776852096408345412394614356", -- LUT(2) = log10 (1.07) = 0.029383777685209640834541239461435646
--		x"0030294705536180071693257673841859", -- LUT(3) = log10 (1.007) = 0.0030294705536180071693257673841859106
--		x"0003038997848124918105176677363847", -- LUT(4) = log10 (1.0007) = 0.00030389978481249181051766773638472442
--		x"0000303995497613986940262206790232", -- LUT(5) = log10 (1.00007) = 0.000030399549761398694026220679023281926
--		x"0000030400507331576102389685938385", -- LUT(6) = log10 (1.000007) = 0.0000030400507331576102389685938385813937
--		x"0000003040060309301778673687882288", -- LUT(7) = log10 (1.0000007) = 3.0400603093017786736878822882945671E-7
--		x"0000000304006126692061969269452039", -- LUT(8) = log10 (1.00000007) = 3.0400612669206196926945203998207159E-8
--		x"0000000030400613626825480365825681", -- LUT(9) = log10 (1.000000007) = 3.0400613626825480365825681585501081E-9
--		x"0000000003040061372258741313391478", -- LUT(10) = log10 (1.0000000007) = 3.0400613722587413133914788120530024E-10
--		x"0000000000304006137321636064549657", -- LUT(11) = log10 (1.00000000007) = 3.0400613732163606454965711682178755E-11
--		x"0000000000030400613733121225787513", -- LUT(12) = log10 (1.000000000007) = 3.0400613733121225787513224169745469E-12
--		x"0000000000003040061373321698772077", -- LUT(13) = log10 (1.0000000000007) = 3.0400613733216987720772399619818480E-13
--		x"0000000000000304006137332265639140", -- LUT(14) = log10 (1.00000000000007) = 3.0400613733226563914098361406838946E-14
--		x"0000000000000030400613733227521533", -- LUT(15) = log10 (1.000000000000007) = 3.0400613733227521533430958027961125E-15
--		x"0000000000000003040061373322761729", -- LUT(16) = log10 (1.0000000000000007) = 3.0400613733227617295364217694497544E-16
--		x"0000000000000000304006137332276268", -- LUT(17) = log10 (1.00000000000000007) = 3.0400613733227626871557543661195428E-17
--		x"0000000000000000030400613733227627", -- LUT(18) = log10 (1.000000000000000007) = 3.0400613733227627829176876257865658E-18
--		x"0000000000000000003040061373322762", -- LUT(19) = log10 (1.0000000000000000007) = 3.0400613733227627924938809517532686E-19
--		x"0000000000000000000304006137332276", -- LUT(20) = log10 (1.00000000000000000007) = 3.0400613733227627934515002843499389E-20
--		x"0000000000000000000030400613733227", -- LUT(21) = log10 (1.000000000000000000007) = 3.0400613733227627935472622176096059E-21
--		x"0000000000000000000003040061373322", -- LUT(22) = log10 (1.0000000000000000000007) = 3.0400613733227627935568384109355726E-22
--		x"0000000000000000000000304006137332", -- LUT(23) = log10 (1.00000000000000000000007) = 3.0400613733227627935577960302681693E-23
--		x"0000000000000000000000030400613733", -- LUT(24) = log10 (1.000000000000000000000007) = 3.0400613733227627935578917922014289E-24
--		x"0000000000000000000000003040061373", -- LUT(25) = log10 (1.0000000000000000000000007) = 3.0400613733227627935579013683947549E-25
--		x"0000000000000000000000000304006137", -- LUT(26) = log10 (1.00000000000000000000000007) = 3.0400613733227627935579023260140875E-26
--		x"0000000000000000000000000030400613", -- LUT(27) = log10 (1.000000000000000000000000007) = 3.0400613733227627935579024217760208E-27
--		x"0000000000000000000000000003040061", -- LUT(28) = log10 (1.0000000000000000000000000007) = 3.0400613733227627935579024313522141E-28
--		x"0000000000000000000000000000304006", -- LUT(29) = log10 (1.00000000000000000000000000007) = 3.0400613733227627935579024323098334E-29
--		x"0000000000000000000000000000030400", -- LUT(30) = log10 (1.000000000000000000000000000007) = 3.0400613733227627935579024324055954E-30
--		x"0000000000000000000000000000003040", -- LUT(31) = log10 (1.0000000000000000000000000000007) = 3.0400613733227627935579024324151716E-31
--		x"0000000000000000000000000000000304", -- LUT(32) = log10 (1.00000000000000000000000000000007) = 3.0400613733227627935579024324161292E-32
--		x"0000000000000000000000000000000030"); -- LUT(33) = log10 (1.000000000000000000000000000000007) = 3.0400613733227627935579024324162249E-33
--
--signal lut_Log10ShN2: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"2552725051033060698037947012347236", -- LUT(1) = log10 (1.8) = 0.25527250510330606980379470123472365
--		x"0334237554869497023125614992143319", -- LUT(2) = log10 (1.08) = 0.033423755486949702312561499214331981
--		x"0034605321095064861572276440008389", -- LUT(3) = log10 (1.008) = 0.0034605321095064861572276440008389190
--		x"0003472966853635406877056930035570", -- LUT(4) = log10 (1.0008) = 0.00034729668536354068770569300355701318
--		x"0000347421688840332004935023775335", -- LUT(5) = log10 (1.00008) = 0.000034742168884033200493502377533561921
--		x"0000034743419578767128640139981982", -- LUT(6) = log10 (1.000008) = 0.0000034743419578767128640139981982054723
--		x"0000003474354465484413726274247152", -- LUT(7) = log10 (1.0000008) = 3.4743544654844137262742471526562701E-7
--		x"0000000347435571625178782412715960", -- LUT(8) = log10 (1.00000008) = 3.4743557162517878241271596009484382E-8
--		x"0000000034743558413285912744245639", -- LUT(9) = log10 (1.000000008) = 3.4743558413285912744245639999341472E-9
--		x"0000000003474355853836272279859821", -- LUT(10) = log10 (1.0000000008) = 3.4743558538362722798598214181860604E-10
--		x"0000000000347435585508704038700740", -- LUT(11) = log10 (1.00000000008) = 3.4743558550870403870074027256418502E-11
--		x"0000000000034743558552121171977882", -- LUT(12) = log10 (1.000000000008) = 3.4743558552121171977882014124395822E-12
--		x"0000000000003474355855224624878866", -- LUT(13) = log10 (1.0000000000008) = 3.4743558552246248788669416866802728E-13
--		x"0000000000000347435585522587564697", -- LUT(14) = log10 (1.00000000000008) = 3.4743558552258756469748223181599515E-14
--		x"0000000000000034743558552260007237", -- LUT(15) = log10 (1.000000000000008) = 3.4743558552260007237856104473484754E-15
--		x"0000000000000003474355855226013231", -- LUT(16) = log10 (1.0000000000000008) = 3.4743558552260132314666892609277334E-16
--		x"0000000000000000347435585522601448", -- LUT(17) = log10 (1.00000000000000008) = 3.4743558552260144822347971422922632E-17
--		x"0000000000000000034743558552260146", -- LUT(18) = log10 (1.000000000000000008) = 3.4743558552260146073116079304287822E-18
--		x"0000000000000000003474355855226014", -- LUT(19) = log10 (1.0000000000000000008) = 3.4743558552260146198192890092424348E-19
--		x"0000000000000000000347435585522601", -- LUT(20) = log10 (1.00000000000000000008) = 3.4743558552260146210700571171238001E-20
--		x"0000000000000000000034743558552260", -- LUT(21) = log10 (1.000000000000000000008) = 3.4743558552260146211951339279119366E-21
--		x"0000000000000000000003474355855226", -- LUT(22) = log10 (1.0000000000000000000008) = 3.4743558552260146212076416089907503E-22
--		x"0000000000000000000000347435585522", -- LUT(23) = log10 (1.00000000000000000000008) = 3.4743558552260146212088923770986316E-23
--		x"0000000000000000000000034743558552", -- LUT(24) = log10 (1.000000000000000000000008) = 3.4743558552260146212090174539094198E-24
--		x"0000000000000000000000003474355855", -- LUT(25) = log10 (1.0000000000000000000000008) = 3.4743558552260146212090299615904986E-25
--		x"0000000000000000000000000347435585", -- LUT(26) = log10 (1.00000000000000000000000008) = 3.4743558552260146212090312123586064E-26
--		x"0000000000000000000000000034743558", -- LUT(27) = log10 (1.000000000000000000000000008) = 3.4743558552260146212090313374354172E-27
--		x"0000000000000000000000000003474355", -- LUT(28) = log10 (1.0000000000000000000000000008) = 3.4743558552260146212090313499430983E-28
--		x"0000000000000000000000000000347435", -- LUT(29) = log10 (1.00000000000000000000000000008) = 3.4743558552260146212090313511938664E-29
--		x"0000000000000000000000000000034743", -- LUT(30) = log10 (1.000000000000000000000000000008) = 3.4743558552260146212090313513189432E-30
--		x"0000000000000000000000000000003474", -- LUT(31) = log10 (1.0000000000000000000000000000008) = 3.4743558552260146212090313513314509E-31
--		x"0000000000000000000000000000000347", -- LUT(32) = log10 (1.00000000000000000000000000000008) = 3.4743558552260146212090313513327017E-32
--		x"0000000000000000000000000000000034"); -- LUT(33) = log10 (1.000000000000000000000000000000008) = 3.4743558552260146212090313513328268E-33
--
--signal lut_Log10ShN1: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"2787536009528289615363334757569293", -- LUT(1) = log10 (1.9) = 0.27875360095282896153633347575692932
--		x"0374264979406236352005133076138752", -- LUT(2) = log10 (1.09) = 0.037426497940623635200513307613875287
--		x"0038911662369105217152813165095588", -- LUT(3) = log10 (1.009) = 0.0038911662369105217152813165095588655
--		x"0003906892499101310288642232545687", -- LUT(4) = log10 (1.0009) = 0.00039068924991013102886422325456872771
--		x"0000390847445841673924188050248845", -- LUT(5) = log10 (1.00009) = 0.000039084744584167392418805024884522862
--		x"0000039086327483082822139172355443", -- LUT(6) = log10 (1.000009) = 0.0000039086327483082822139172355443443391
--		x"0000003908648578237670075568932174", -- LUT(7) = log10 (1.0000009) = 3.9086485782376700755689321740694201E-7
--		x"0000000390865016124001183139836796", -- LUT(8) = log10 (1.00000009) = 3.9086501612400118313983679690889930E-8
--		x"0000000039086503195403400373120196", -- LUT(9) = log10 (1.000000009) = 3.9086503195403400373120196405173998E-9
--		x"0000000003908650335370373798207325", -- LUT(10) = log10 (1.0000000009) = 3.9086503353703737982073259585749240E-10
--		x"0000000000390865033695337718369989", -- LUT(11) = log10 (1.00000000009) = 3.9086503369533771836998966359602752E-11
--		x"0000000000039086503371116775223431", -- LUT(12) = log10 (1.000000000009) = 3.9086503371116775223431841047886768E-12
--		x"0000000000003908650337127507556208", -- LUT(13) = log10 (1.0000000000009) = 3.9086503371275075562084531556830497E-13
--		x"0000000000000390865033712909055959", -- LUT(14) = log10 (1.00000000000009) = 3.9086503371290905595949894638126029E-14
--		x"0000000000000039086503371292488599", -- LUT(15) = log10 (1.000000000000009) = 3.9086503371292488599336431886559594E-15
--		x"0000000000000003908650337129264689", -- LUT(16) = log10 (1.0000000000000009) = 3.9086503371292646899675085620805991E-16
--		x"0000000000000000390865033712926627", -- LUT(17) = log10 (1.00000000000000009) = 3.9086503371292662729708950994324661E-17
--		x"0000000000000000039086503371292664", -- LUT(18) = log10 (1.000000000000000009) = 3.9086503371292664312712337531677468E-18
--		x"0000000000000000003908650337129266", -- LUT(19) = log10 (1.0000000000000000009) = 3.9086503371292664471012676185412758E-19
--		x"0000000000000000000390865033712926", -- LUT(20) = log10 (1.00000000000000000009) = 3.9086503371292664486842710050786288E-20
--		x"0000000000000000000039086503371292", -- LUT(21) = log10 (1.000000000000000000009) = 3.9086503371292664488425713437323640E-21
--		x"0000000000000000000003908650337129", -- LUT(22) = log10 (1.0000000000000000000009) = 3.9086503371292664488584013775977376E-22
--		x"0000000000000000000000390865033712", -- LUT(23) = log10 (1.00000000000000000000009) = 3.9086503371292664488599843809842749E-23
--		x"0000000000000000000000039086503371", -- LUT(24) = log10 (1.000000000000000000000009) = 3.9086503371292664488601426813229287E-24
--		x"0000000000000000000000003908650337", -- LUT(25) = log10 (1.0000000000000000000000009) = 3.9086503371292664488601585113567940E-25
--		x"0000000000000000000000000390865033", -- LUT(26) = log10 (1.00000000000000000000000009) = 3.9086503371292664488601600943601806E-26
--		x"0000000000000000000000000039086503", -- LUT(27) = log10 (1.000000000000000000000000009) = 3.9086503371292664488601602526605192E-27
--		x"0000000000000000000000000003908650", -- LUT(28) = log10 (1.0000000000000000000000000009) = 3.9086503371292664488601602684905531E-28
--		x"0000000000000000000000000000390865", -- LUT(29) = log10 (1.00000000000000000000000000009) = 3.9086503371292664488601602700735565E-29
--		x"0000000000000000000000000000039086", -- LUT(30) = log10 (1.000000000000000000000000000009) = 3.9086503371292664488601602702318568E-30
--		x"0000000000000000000000000000003908", -- LUT(31) = log10 (1.0000000000000000000000000000009) = 3.9086503371292664488601602702476868E-31
--		x"0000000000000000000000000000000390", -- LUT(32) = log10 (1.00000000000000000000000000000009) = 3.9086503371292664488601602702492699E-32
--		x"0000000000000000000000000000000039"); -- LUT(33) = log10 (1.000000000000000000000000000000009) = 3.9086503371292664488601602702494282E-33
--
--signal lut_Log10ShN0: mlut_LogShN := (
--		x"0000000000000000000000000000000000", -- LUT(0), No usada
--		x"3010299956639811952137388947244930", -- LUT(1) = log10 (2.0) = 0.30102999566398119521373889472449303
--		x"0413926851582250407501999712430242", -- LUT(2) = log10 (1.10) = 0.041392685158225040750199971243024242
--		x"0043213737826425742751881782229379", -- LUT(3) = log10 (1.010) = 0.0043213737826425742751881782229379132
--		x"0004340774793186406689213877779888", -- LUT(4) = log10 (1.0010) = 0.00043407747931864066892138777798886602
--		x"0000434272768626696373135275850982", -- LUT(5) = log10 (1.00010) = 0.000043427276862669637313527585098268131
--		x"0000043429231044531868554934716343", -- LUT(6) = log10 (1.000010) = 0.0000043429231044531868554934716343971840
--		x"0000004342942647561556407439426436", -- LUT(7) = log10 (1.0000010) = 4.3429426475615564074394264367770704E-7
--		x"0000000434294460188529180136701973", -- LUT(8) = log10 (1.00000010) = 4.3429446018852918013670197358779472E-8
--		x"0000000043429447973177943261135240", -- LUT(9) = log10 (1.000000010) = 4.3429447973177943261135240219573514E-9
--		x"0000000004342944816861045868442678", -- LUT(10) = log10 (1.0000000010) = 4.3429448168610458684426783228355094E-10
--		x"0000000000434294481881537103557413", -- LUT(11) = log10 (1.00000000010) = 4.3429448188153710355741397580695090E-11
--		x"0000000000043429448190108035524162", -- LUT(12) = log10 (1.000000000010) = 4.3429448190108035524162713626107944E-12
--		x"0000000000004342944819030346804101", -- LUT(13) = log10 (1.0000000000010) = 4.3429448190303468041017743776760682E-13
--		x"0000000000000434294481903230112927", -- LUT(14) = log10 (1.00000000000010) = 4.3429448190323011292703375777287080E-14
--		x"0000000000000043429448190324965617", -- LUT(15) = log10 (1.000000000000010) = 4.3429448190324965617871940267194331E-15
--		x"0000000000000004342944819032516105", -- LUT(16) = log10 (1.0000000000000010) = 4.3429448190325161050388796729083602E-16
--		x"0000000000000000434294481903251805", -- LUT(17) = log10 (1.00000000000000010) = 4.3429448190325180593640482375401515E-17
--		x"0000000000000000043429448190325182", -- LUT(18) = log10 (1.000000000000000010) = 4.3429448190325182547965650940034596E-18
--		x"0000000000000000004342944819032518", -- LUT(19) = log10 (1.0000000000000000010) = 4.3429448190325182743398167796497917E-19
--		x"0000000000000000000434294481903251", -- LUT(20) = log10 (1.00000000000000000010) = 4.3429448190325182762941419482144249E-20
--		x"0000000000000000000043429448190325", -- LUT(21) = log10 (1.000000000000000000010) = 4.3429448190325182764895744650708882E-21
--		x"0000000000000000000004342944819032", -- LUT(22) = log10 (1.0000000000000000000010) = 4.3429448190325182765091177167565346E-22
--		x"0000000000000000000000434294481903", -- LUT(23) = log10 (1.00000000000000000000010) = 4.3429448190325182765110720419250992E-23
--		x"0000000000000000000000043429448190", -- LUT(24) = log10 (1.000000000000000000000010) = 4.3429448190325182765112674744419557E-24
--		x"0000000000000000000000004342944819", -- LUT(25) = log10 (1.0000000000000000000000010) = 4.3429448190325182765112870176936413E-25
--		x"0000000000000000000000000434294481", -- LUT(26) = log10 (1.00000000000000000000000010) = 4.3429448190325182765112889720188099E-26
--		x"0000000000000000000000000043429448", -- LUT(27) = log10 (1.000000000000000000000000010) = 4.3429448190325182765112891674513267E-27
--		x"0000000000000000000000000004342944", -- LUT(28) = log10 (1.0000000000000000000000000010) = 4.3429448190325182765112891869945784E-28
--		x"0000000000000000000000000000434294", -- LUT(29) = log10 (1.00000000000000000000000000010) = 4.3429448190325182765112891889489036E-29
--		x"0000000000000000000000000000043429", -- LUT(30) = log10 (1.000000000000000000000000000010) = 4.3429448190325182765112891891443361E-30
--		x"0000000000000000000000000000004342", -- LUT(31) = log10 (1.0000000000000000000000000000010) = 4.3429448190325182765112891891638794E-31
--		x"0000000000000000000000000000000434", -- LUT(32) = log10 (1.00000000000000000000000000000010) = 4.3429448190325182765112891891658337E-32
--		x"0000000000000000000000000000000043"); -- LUT(33) = log10 (1.000000000000000000000000000000010) = 4.3429448190325182765112891891660291E-33
--
--

-- ====== FIN declaraci�n
-- declaracion de meomria de ln para la parte de x<1

type mem_LogSh_P is array (0 to 9) of STD_LOGIC_VECTOR (4*P-1 downto 0); 
type mem_LogSh_N is array (0 to 9) of STD_LOGIC_VECTOR (4*P-1 downto 0); 

signal vlog_ShP: mem_LogSh_P;
signal vlog_ShN: mem_LogSh_N;

signal log_ShPN, log_Sh0: std_logic_vector(4*P downto 0);

begin

	vlog_ShP(0) <= (others => '0');
	vlog_ShP(1) <= lut_Log10ShP1(conv_integer(step));
	vlog_ShP(2) <= lut_Log10ShP2(conv_integer(step));
	vlog_ShP(3) <= lut_Log10ShP3(conv_integer(step));
	vlog_ShP(4) <= lut_Log10ShP4(conv_integer(step));
	vlog_ShP(5) <= lut_Log10ShP5(conv_integer(step));
	vlog_ShP(6) <= lut_Log10ShP6(conv_integer(step));
	vlog_ShP(7) <= lut_Log10ShP7(conv_integer(step));
	vlog_ShP(8) <= lut_Log10ShP8(conv_integer(step));
	vlog_ShP(9) <= lut_Log10ShP9(conv_integer(step));

	vlog_ShN(0) <= lut_Log10ShN0(conv_integer(step));
	vlog_ShN(1) <= lut_Log10ShN1(conv_integer(step));
	vlog_ShN(2) <= lut_Log10ShN2(conv_integer(step));
	vlog_ShN(3) <= lut_Log10ShN3(conv_integer(step));
	vlog_ShN(4) <= lut_Log10ShN4(conv_integer(step));
	vlog_ShN(5) <= lut_Log10ShN5(conv_integer(step));
	vlog_ShN(6) <= lut_Log10ShN6(conv_integer(step));
	vlog_ShN(7) <= lut_Log10ShN7(conv_integer(step));
	vlog_ShN(8) <= lut_Log10ShN8(conv_integer(step));
	vlog_ShN(9) <= lut_Log10ShN9(conv_integer(step));

	
	log_ShPN(4*P-1 downto 0) <= vlog_ShP(conv_integer(d)) when (x_greater_1='1') else vlog_ShN(conv_integer(d));
	log_ShPN(4*P) <= x_greater_1;
	
	log_Sh0(4*P) <= '0';
	log_Sh0(4*P-1 downto 0) <= lut_Log(conv_integer(d));
	
	
	log <= log_Sh0 when (step_eq_0='1') else log_ShPN;	


end Behavioral;

