

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.my_package.all;

Library UNISIM;
use UNISIM.vcomponents.all;

entity Lutb_log_pf34_bopt is
	generic (P: integer:=34);
    port ( 
 			step : in std_logic_vector(log2sup(P+2)-1 downto 0);
			offset_step : in std_logic_vector(log2sup(P+1)-1 downto 0);
			true_step: in std_logic_vector(log2sup(2*P+1)-1 downto 0);
           d : in  STD_LOGIC_VECTOR (3 downto 0);-- corresponde a xi
			  x_greater_1: in std_logic; -- indica si x es mayor a uno
           log : out  STD_LOGIC_VECTOR (4*P+8 downto 0)); -- en SVA, por eso un bit m�s
end Lutb_log_pf34_bopt;


architecture Behavioral of Lutb_log_pf34_bopt is


-- == Comienzo declaraci�n

	
-- ====== Comienzo declaraci�n
-- declaracion de meomria de log para la parte de x>1
-- Precisi�n 35

type mlut_LogShP is array (0 to P+2) of std_logic_vector (8*P+7 downto 0);

signal lut_LogShP1: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"0457574905606750002560000000000013815997422716186082703402687193895411", -- LUT(1) = log (0.9) = -0.045757490560675125409944193489769381599742271618608270340268719389541694
		x"0043648054024500000512000000000001398930400811521551757437297007097882", -- LUT(2) = log (0.99) = -0.0043648054024500846597442222467451398930400811521551757437297007097886622
		x"0004345117740176900051200000000000144166407172615998588927231682907273", -- LUT(3) = log (0.999) = -0.00043451177401769130646560069552462441664071726159985889272316829072711623
		x"0000434316198075100005120000000000016737507259457025843379110637613400", -- LUT(4) = log (0.9999) = -0.000043431619807510384556044023807226673750725945702584337911063761340651830
		x"0000043429665339013000512000000000001412005380734464616369437218737994", -- LUT(5) = log (0.99999) = -0.0000043429665339013793521486464083130412005380734464616369437218737997944893
		x"0000004342946990506300025600000000000166369420841130859913582208951675", -- LUT(6) = log (0.999999) = -4.3429469905063754421291753575839663694208411308599135822089516755246202E-7
		x"0000000434294503617970000000000000000018235206516193204036885358451336", -- LUT(7) = log (0.9999999) = -4.3429450361797737046210188594163823520651619320403688535845133809805530E-8
		x"0000000043429448407472000000000000000001527631698100535646646595497557", -- LUT(8) = log (0.99999999) = -4.3429448407472425164387089585426527631698100535646646595497558928195276E-9
		x"0000000004342944821203900076800000000000171048657477066222151054197137", -- LUT(9) = log (0.999999999) = -4.3429448212039906874751966015182710486574770662221510541971382935403065E-10
		x"0000000000434294481924960000000000000000010941286215521827993337769377", -- LUT(10) = log (0.9999999999) = -4.3429448192496655174773915857228094128621552182799333776937050946833309E-11
		x"0000000000043429448190542000000000000000001094385685554552731498124217", -- LUT(11) = log (0.99999999999) = -4.3429448190542330006065965453759094385685554552731498124218688838194169E-12
		x"0000000000004342944819034600025600000000000179479463714791970198859619", -- LUT(12) = log (0.999999999999) = -4.3429448190346897489208068959525794794637147919701988596154600039168562E-13
		x"0000000000000434294481903270000000000000000015911751290835182020170668", -- LUT(13) = log (0.9999999999999) = -4.3429448190327354237522408295563591175129083518202017066289666110431659E-14
		x"0000000000000043429448190325000768000000000001982066910009165773614457", -- LUT(14) = log (0.99999999999999) = -4.3429448190325399912353843519021982066910009165773614454386180598787803E-15
		x"0000000000000004342944819032500025600000000000136726861575481573317106", -- LUT(15) = log (0.999999999999999) = -4.3429448190325204479836987054266367268615754815733171009507526379825778E-16
		x"0000000000000000434294481903250007680000000000017912499115962473454755", -- LUT(16) = log (0.9999999999999999) = -4.3429448190325184936585301407919791249911596247345475821784294166506594E-17
		x"0000000000000000043429448190325000768000000000001423502652433049508634", -- LUT(17) = log (0.99999999999999999) = -4.3429448190325182982260132843286423502652433049508634119768991855065800E-18
		x"0000000000000000004342944819032500076800000000000109962647262925630533", -- LUT(18) = log (0.999999999999999999) = -4.3429448190325182786827615986823099626472629256305304992060221284904592E-19
		x"0000000000000000000434294481903250005120000000000017673678401100022502", -- LUT(19) = log (0.9999999999999999999) = -4.3429448190325182767284364301176767367840110002250765965478597013957914E-20
		x"0000000000000000000043429448190325000512000000000001134143266712688094", -- LUT(20) = log (0.99999999999999999999) = -4.3429448190325182765330039132612134143266712688097969992018091439913401E-21
		x"0000000000000000000004342944819032500051200000000000167082082227150272", -- LUT(21) = log (0.999999999999999999999) = -4.3429448190325182765134606615755670820822271502795216973954353215364641E-22
		x"0000000000000000000000434294481903250005120000000000010244885779563690", -- LUT(22) = log (0.9999999999999999999999) = -4.3429448190325182765115063364070024488577956369726066937940792852002647E-23
		x"0000000000000000000000043429448190325000512000000000001459855353526140", -- LUT(23) = log (0.99999999999999999999999) = -4.3429448190325182765113109038901459855353526146273763186997364940593141E-24
		x"0000000000000000000000004342944819032500051200000000000160339203108315", -- LUT(24) = log (0.999999999999999999999999) = -4.3429448190325182765112913606384603392031083136827078924429601430691793E-25
		x"0000000000000000000000000434294481903250005120000000000019177456988387", -- LUT(25) = log (0.9999999999999999999999999) = -4.3429448190325182765112894063132917745698838836011395959298090872514044E-26
		x"0000000000000000000000000043429448190325000512000000000001749181065618", -- LUT(26) = log (0.99999999999999999999999999) = -4.3429448190325182765112892108807749181065614405931117517396192474624393E-27
		x"0000000000000000000000000004342944819032500051200000000000123232460226", -- LUT(27) = log (0.999999999999999999999999999) = -4.3429448190325182765112891913375232324602291962923102571752115161414709E-28
		x"0000000000000000000000000000434294481903250005120000000000019806389551", -- LUT(28) = log (0.9999999999999999999999999999) = -4.3429448190325182765112891893831980638955959718622301206173168555359534E-29
		x"0000000000000000000000000000043429448190325000512000000000001655470390", -- LUT(29) = log (0.99999999999999999999999999999) = -4.3429448190325182765112891891877655470391326494192221070905128506006674E-30
		x"0000000000000000000000000000004342944819032500051200000000000122295350", -- LUT(30) = log (0.999999999999999999999999999999) = -4.3429448190325182765112891891682222953534863171749213057391223047183915E-31
		x"0000000000000000000000000000000434294481903250005120000000000016797010", -- LUT(31) = log (0.9999999999999999999999999999999) = -4.3429448190325182765112891891662679701849216839504912256039961486762764E-32
		x"0000000000000000000000000000000043429448190325000512000000000001725379", -- LUT(32) = log (0.99999999999999999999999999999999) = -4.3429448190325182765112891891660725376680652206280482175904836620575260E-33
		x"0000000000000000000000000000000004342944819032500051200000000000152998", -- LUT(33) = log (0.999999999999999999999999999999999) = -4.3429448190325182765112891891660529944163795742958039167891324146855056E-34
		x"0000000000000000000000000000000000434294481903250005120000000000015106", -- LUT(34) = log (0.9999999999999999999999999999999999) = -4.3429448190325182765112891891660510400912110096625794867089972899612021E-35
		x"0000000000000000000000000000000000043429448190325000512000000000001506", -- LUT(35) = log (0.99999999999999999999999999999999999) = -4.3429448190325182765112891891660508446586941531992570437009837774889008E-36
		x"0000000000000000000000000000000000004342944819032500051200000000000150"); -- LUT(36) = log (0.999999999999999999999999999999999999) = -4.3429448190325182765112891891660508446586941531992570437009837774889008E-37
		
		
signal lut_LogShP2: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"0969100130080560002560000000000019196954303556136743760687176166186751", -- LUT(1) = log (0.8) = -0.096910013008056414358783315826520919695430355613674376068717616618675432
		x"0087739243075051000512000000000001862646653258899606456823026314363840", -- LUT(2) = log (0.98) = -0.0087739243075051433618285880902345862646653258899606456823026314363849309
		x"0008694587126288900000000000000000159155412287720410179678859386076842", -- LUT(3) = log (0.998) = -0.00086945871262889062035606924211850591554122877204101796788593860768405165
		x"0000868675834285800005120000000000010461114135647978614370065895055903", -- LUT(4) = log (0.9998) = -0.000086867583428580794567691758055002046111413564797861437006589505590219929
		x"0000086859764981195000768000000000001715047748208277059658891945595234", -- LUT(5) = log (0.99998) = -0.0000086859764981195531938540093755639715047748208277059658891945595237130912
		x"0000008685898323966200000000000000000149820806489190672136582683282185", -- LUT(6) = log (0.999998) = -8.6858983239662558216150251873377498208064891906721365826832821874594828E-7
		x"0000000868589050665410005120000000000019500067753276394381042537364556", -- LUT(7) = log (0.9999998) = -8.6858905066541161714054463297995950006775327639438104253736455025570042E-8
		x"0000000086858897249239000768000000000001799107655636201124538571299427", -- LUT(8) = log (0.99999998) = -8.6858897249239340917915796890089799107655636201124538571299422704876659E-9
		x"0000000008685889646750900000000000000000174732175066260582092174976828", -- LUT(9) = log (0.999999998) = -8.6858896467509262026688011328131747321750662605820921749768244506891645E-10
		x"0000000000868588963893360000000000000000019841704036088349724257174269", -- LUT(10) = log (0.9999999998) = -8.6858896389336255169448938954925984170403608834972425717426556412643150E-11
		x"0000000000086858896381518000256000000000001534729909405510042294715397", -- LUT(11) = log (0.99999999998) = -8.6858896381518954494043868624807534729909405510042294715396615365288934E-12
		x"0000000000008685889638073700025600000000000108328353455523981591658095", -- LUT(12) = log (0.999999999998) = -8.6858896380737224426606549960713083283534555239815916580943547102716821E-13
		x"0000000000000868588963806590002560000000000016574461029914581509801334", -- LUT(13) = log (0.9999999999998) = -8.6858896380659051419863849977992657446102991458150980133194342796536654E-14
		x"0000000000000086858896380651000000000000000001504900804123492720767823", -- LUT(14) = log (0.99999999999998) = -8.6858896380651234119189590298557504900804123492720767824855711296570837E-15
		x"0000000000000008685889638065000025600000000000135854650405180950786592", -- LUT(15) = log (0.999999999999998) = -8.6858896380650452389122164433802358546504051809507865908637354397351311E-16
		x"0000000000000000868588963806500000000000000000017276000761881645490791", -- LUT(16) = log (0.9999999999999998) = -8.6858896380650374216115421848358727600076188164549079914042617745579002E-17
		x"0000000000000000086858896380650000256000000000001683342323423080659058", -- LUT(17) = log (0.99999999999999998) = -8.6858896380650366398814747589824683342323423080659055559582033984042097E-18
		x"0000000000000000008685889638065000051200000000000138210491704678492149", -- LUT(18) = log (0.999999999999999998) = -8.6858896380650365617084680163971382104917046784921483895788995599634996E-19
		x"0000000000000000000868588963806500005120000000000010530130600981574749", -- LUT(19) = log (0.9999999999999999998) = -8.6858896380650365538911673421386053013060098157474086409355424992451842E-20
		x"0000000000000000000086858896380650000512000000000001520114193240184752", -- LUT(20) = log (0.99999999999999999998) = -8.6858896380650365531094372747127520114193240184750610102883754467077467E-21
		x"0000000000000000000008685889638065000051200000000000166682440974275630", -- LUT(21) = log (0.999999999999999999998) = -8.6858896380650365530312642679701666824409742756378475106503676509096500E-22
		x"0000000000000000000000868588963806500005120000000000010814954324248973", -- LUT(22) = log (0.9999999999999999999998) = -8.6858896380650365530234469672959081495432424897230263733208184976473171E-23
		x"0000000000000000000000086858896380650000512000000000001822962534703434", -- LUT(23) = log (0.99999999999999999999998) = -8.6858896380650365530226652372284822962534703430152332617142060831214815E-24
		x"0000000000000000000000008685889638065000051200000000000139710924493131", -- LUT(24) = log (0.999999999999999999999998) = -8.6858896380650365530225870642217397109244931386632908405748082666614392E-25
		x"0000000000000000000000000868588963806500005120000000000016545239159548", -- LUT(25) = log (0.9999999999999999999999998) = -8.6858896380650365530225792469210654523915954183312849673610811192653449E-26
		x"0000000000000000000000000086858896380650000512000000000001980265383056", -- LUT(26) = log (0.99999999999999999999999998) = -8.6858896380650365530225784651909980265383056462991162637287105308682345E-27
		x"0000000000000000000000000008685889638065000051200000000000191283952976", -- LUT(27) = log (0.999999999999999999999999998) = -8.6858896380650365530225783870179912839529766690959097122023634932919485E-28
		x"0000000000000000000000000000868588963806500005120000000000019060969445", -- LUT(28) = log (0.9999999999999999999999999998) = -8.6858896380650365530225783792006906096944437713755891602380976897469541E-29
		x"0000000000000000000000000000086858896380650000512000000000001605422680", -- LUT(29) = log (0.99999999999999999999999999998) = -8.6858896380650365530225783784189605422685904816035571060735547983945811E-30
		x"0000000000000000000000000000008685889638065000051200000000000187535520", -- LUT(30) = log (0.999999999999999999999999999998) = -8.6858896380650365530225783783407875355260051526263539006674193461493650E-31
		x"0000000000000000000000000000000868588963806500005120000000000017023485", -- LUT(31) = log (0.9999999999999999999999999999998) = -8.6858896380650365530225783783329702348517466197286335801269089892937436E-32
		x"0000000000000000000000000000000086858896380650000512000000000001885044", -- LUT(32) = log (0.99999999999999999999999999999998) = -8.6858896380650365530225783783321885047843207664388615480728589854918705E-33
		x"0000000000000000000000000000000008685889638065000051200000000000110333", -- LUT(33) = log (0.999999999999999999999999999999998) = -8.6858896380650365530225783783321103317775781811098843448674539954305201E-34
		x"0000000000000000000000000000000000868588963806500005120000000000010252", -- LUT(34) = log (0.9999999999999999999999999999999998) = -8.6858896380650365530225783783321025144769039225769866245469134965275734E-35
		x"0000000000000000000000000000000000086858896380650000512000000000001010",-- LUT(35) = log (0.99999999999999999999999999999999998) = -8.6858896380650365530225783783321017327468364967236968525148594466383106E-36
		x"0000000000000000000000000000000000008685889638065000051200000000000101"); -- LUT(36) = log (0.999999999999999999999999999999999998) = -8.6858896380650365530225783783321017327468364967236968525148594466383106E-37
		
signal lut_LogShP3: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"1549019599857400076800000000000138065164276036760345934963650462817460", -- LUT(1) = log (0.7) = -0.15490195998574316928778374140736380651642760367603459349636504628174656
		x"0132282657337550000000000000000015505741584153611330252812793271104465", -- LUT(2) = log (0.97) = -0.013228265733755148215638188334422550574158415361133025281279327110446007
		x"0013048416883442000000000000000001072908709904374765421762885821898166", -- LUT(3) = log (0.997) = -0.0013048416883442801186282971867276072908709904374765421762885821898161990
		x"0001303078917321900076800000000000136264465448761684742447793109173521", -- LUT(4) = log (0.9997) = -0.00013030789173219118920260206698228362644654487616847424477931091735261198
		x"0000130290298935230005120000000000011753565854852847183588076320064742", -- LUT(5) = log (0.99997) = -0.000013029029893523149576728886383053175356585485284718358807632006474580677
		x"0000013028854000388000000000000000001474550881010749808106119576562593", -- LUT(6) = log (0.999997) = -0.0000013028854000388327067182248185842474550881010749808106119576562592863333
		x"0000001302883641142300025600000000000129920185850985830755130927046624", -- LUT(7) = log (0.9999997) = -1.3028836411423114259288749577915299201858509858307551309270466237554239E-7
		x"0000000130288346525300005120000000000013109211943833944309605220123545", -- LUT(8) = log (0.99999997) = -1.3028834652530075594647615084407310921194383394430960522012354459075184E-8
		x"0000000013028834476640000512000000000001251105156355411854110839466546", -- LUT(9) = log (0.999999997) = -1.3028834476640806554266703271036251105156355411854110839466543011866433E-9
		x"0000000001302883445905100076800000000000110388144916427838485640647607", -- LUT(10) = log (0.9999999997) = -1.3028834459051879998489365825729103881449164278384856406476009112090165E-10
		x"0000000000130288344572920002560000000000013776934258301405790065379628", -- LUT(11) = log (0.99999999997) = -1.3028834457292987346394239540278377693425830140579006537962655572397344E-11
		x"0000000000013028834457117000000000000000001824650792278590035509560719", -- LUT(12) = log (0.999999999997) = -1.3028834457117098081219552986245824650792278590035509560711299122828104E-12
		x"0000000000001302883445709900000000000000000161626198162441558177839670", -- LUT(13) = log (0.9999999999997) = -1.3028834457099509154702432591587616261981624415581778396715478168876874E-13
		x"0000000000000130288344570970002560000000000012458139747770398897751429", -- LUT(14) = log (0.99999999999997) = -1.3028834457097750262050724034729245813974777039889775142941441421236201E-14
		x"0000000000000013028834457097000256000000000001483273004554173771934418", -- LUT(15) = log (0.999999999999997) = -1.3028834457097574372785553213869483273004554173771934419410075283849721E-15
		x"0000000000000001302883445709700076800000000000176776394575822556569796", -- LUT(16) = log (0.9999999999999997) = -1.3028834457097556783859036132131767763945758225565697956832573072255617E-16
		x"0000000000000000130288344570970000000000000000014788204902608158488205", -- LUT(17) = log (0.99999999999999997) = -1.3028834457097555024966384423961478820490260815848820820705121764568845E-17
		x"0000000000000000013028834457097000768000000000001484752219214896649897", -- LUT(18) = log (0.999999999999999997) = -1.3028834457097554849077119253144484752219214896649890263227714044043888E-18
		x"0000000000000000001302883445709700076800000000000178569365285534294764", -- LUT(19) = log (0.9999999999999999997) = -1.3028834457097554831488192736062785693652855342947646498732360680702792E-19
		x"0000000000000000000130288344570970007680000000000016157912788268379593", -- LUT(20) = log (0.99999999999999999997) = -1.3028834457097554829729300084354615791278826837959598536915040252490424E-20
		x"0000000000000000000013028834457097000768000000000001798801076250061962", -- LUT(21) = log (0.999999999999999999997) = -1.3028834457097554829553410819183798801076250061964615504801350049784440E-21
		x"0000000000000000000001302883445709700076800000000000171710205634064511", -- LUT(22) = log (0.9999999999999999999997) = -1.3028834457097554829535821892666717102056340645110155419230583167606028E-22
		x"0000000000000000000000130288344570970007680000000000010089321543531868", -- LUT(23) = log (0.99999999999999999999997) = -1.3028834457097554829534063000015008932154353186032159792849912422488799E-23
		x"0000000000000000000000013028834457097000768000000000001838115164154470", -- LUT(24) = log (0.999999999999999999999997) = -1.3028834457097554829533887110749838115164154474950434734033609407329802E-24
		x"0000000000000000000000001302883445709700076800000000000132103346513460", -- LUT(25) = log (0.9999999999999999999999997) = -1.3028834457097554829533869521823321033465134604190522973190196746407352E-25
		x"0000000000000000000000000130288344570970007680000000000016693252952326", -- LUT(26) = log (0.99999999999999999999999997) = -1.3028834457097554829533867762930669325295232617118014404556237656721041E-26
		x"0000000000000000000000000013028834457097000768000000000001404154478246", -- LUT(27) = log (0.999999999999999999999999997) = -1.3028834457097554829533867587041404154478242418410798373767345569516469E-27
		x"0000000000000000000000000001302883445709700076800000000000147763739656", -- LUT(28) = log (0.9999999999999999999999999997) = -1.3028834457097554829533867569452477637396543398540077118949201399013653E-28
		x"0000000000000000000000000000130288344570970007680000000000015849856881", -- LUT(29) = log (0.99999999999999999999999999997) = -1.3028834457097554829533867567693584985688373496553004996949994432345547E-29
		x"0000000000000000000000000000013028834457097000768000000000001695720512", -- LUT(30) = log (0.999999999999999999999999999997) = -1.3028834457097554829533867567517695720517556506354297784784899810182559E-30
		x"0000000000000000000000000000001302883445709700076800000000000110679403", -- LUT(31) = log (0.9999999999999999999999999999997) = -1.3028834457097554829533867567500106794000474807334427063568738608711298E-31
		x"0000000000000000000000000000000130288344570970007680000000000013479014", -- LUT(32) = log (0.99999999999999999999999999999997) = -1.3028834457097554829533867567498347901348766637432439991447125971171622E-32
		x"0000000000000000000000000000000013028834457097000768000000000001172015", -- LUT(33) = log (0.999999999999999999999999999999997) = -1.3028834457097554829533867567498172012083595820442241284234964742243729E-33
		x"0000000000000000000000000000000001302883445709700076800000000000115446", -- LUT(34) = log (0.9999999999999999999999999999999997) = -1.3028834457097554829533867567498154423157078738743221413513748619699201E-34
		x"0000000000000000000000000000000000130288344570970007680000000000011527", -- LUT(35) = log (0.99999999999999999999999999999999997) = -1.3028834457097554829533867567498152664264427030573319426441627007448230E-35
		x"0000000000000000000000000000000000013028834457097000768000000000001152"); -- LUT(36) = log (0.999999999999999999999999999999999997) = -1.3028834457097554829533867567498152664264427030573319426441627007448230E-36

signal lut_LogShP4: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2218487496163500051200000000000116640316812543471955938597068985676624", -- LUT(1) = log (0.6) = -0.22184874961635636749123320202039166403168125434719559385970689856766266
		x"0177287669604310005120000000000015569589217284987614286179970540592293", -- LUT(2) = log (0.96) = -0.017728766960431586636277623122419556958921728498761428617997054059229901
		x"0017406615763012000256000000000001902618537148044565990199086088722734", -- LUT(3) = log (0.996) = -0.0017406615763012684447339552686373902618537148044565990199086088722732495
		x"0001737525455875800025600000000000102887792018121098421616410476593535", -- LUT(4) = log (0.9996) = -0.00017375254558758231289189578228922028877920181210984216164104765935352661
		x"0000173721267209800005120000000000013552980931273778947464509562750640", -- LUT(5) = log (0.99996) = -0.000017372126720980822612139715542103355298093127377894746450956275064054716
		x"0000017371814019781000000000000000001858840817879783829206293095090830", -- LUT(6) = log (0.999996) = -0.0000017371814019781275133613420426354858840817879783829206293095090832439158
		x"0000001737178275048600076800000000000149774430638706066456610440727460", -- LUT(7) = log (0.9999996) = -1.7371782750486854827232453460289497744306387060664566104407274666934488E-7
		x"0000000173717796235650007680000000000019740815991033183220174782333236", -- LUT(8) = log (0.99999996) = -1.7371779623565667893595844095416974081599103318322017478233323717411505E-8
		x"0000000017371779310873000512000000000001709344861394450606765092320525", -- LUT(9) = log (0.999999996) = -1.7371779310873631750954792719396709344861394450606765092320521429130853E-9
		x"0000000001737177927960400076800000000000112034393815393047741918561989", -- LUT(10) = log (0.9999999996) = -1.7371779279604428962197666272878120343938153930477419185619869553857738E-10
		x"0000000000173717792764770005120000000000016537477008153571064208885607", -- LUT(11) = log (0.99999999996) = -1.7371779276477508691577023167732653747700815357106420888560601627474442E-11
		x"0000000000017371779276164000512000000000001766576960909298536854743124", -- LUT(12) = log (0.999999999996) = -1.7371779276164816664597509552365766576960909298536854743123333423271548E-12
		x"0000000000001737177927613300025600000000000130705034239386363154828923", -- LUT(13) = log (0.9999999999996) = -1.7371779276133547461900383697780307050342393863631548289255372544272547E-13
		x"0000000000000173717792761300005120000000000012731421806637879049998552", -- LUT(14) = log (0.99999999999996) = -1.7371779276130420541630679367391273142180663787904999855801083727388281E-14
		x"0000000000000017371779276130000768000000000001064871562087561733955451", -- LUT(15) = log (0.999999999999996) = -1.7371779276130107849603709016903064871562087561733955450456217169337459E-15
		x"0000000000000001737177927613000051200000000000175099570195850249759183", -- LUT(16) = log (0.9999999999999996) = -1.7371779276130076580401011982679750995701958502497591876532634438782909E-16
		x"0000000000000000173717792761300002560000000000016746776279626348033294", -- LUT(17) = log (0.99999999999999996) = -1.7371779276130073453480742279265674677627962634803329652647777604988186E-17
		x"0000000000000000017371779276130000000000000000001349596515683218168795", -- LUT(18) = log (0.999999999999999996) = -1.7371779276130073140788715308924349596515683218168792738319216244551499E-18
		x"0000000000000000001737177927613000000000000000000121791391140647820646", -- LUT(19) = log (0.9999999999999999996) = -1.7371779276130073109519512611890217913911406478206440535533684201837424E-19
		x"0000000000000000000173717792761300000000000000000018047539060483162277", -- LUT(20) = log (0.99999999999999999996) = -1.7371779276130073106392592342186804753906048316227216082737170963349492E-20
		x"0000000000000000000017371779276130000000000000000001463437988063195148", -- LUT(21) = log (0.999999999999999999996) = -1.7371779276130073106079900315216463437988063195149463744884935605883383E-21
		x"0000000000000000000001737177927613000000000000000000142930639709018999", -- LUT(22) = log (0.9999999999999999999996) = -1.7371779276130073106048631112519429306397090189992890212173738825367324E-22
		x"0000000000000000000000173717792761300000000000000000017258932380011440", -- LUT(23) = log (0.99999999999999999999996) = -1.7371779276130073106045504192249725893238001144546744875913359167463590E-23
		x"0000000000000000000000017371779276130000000000000000001755551922092320", -- LUT(24) = log (0.999999999999999999999996) = -1.7371779276130073106045191500222755551922092322552825462457428601627291E-24
		x"0000000000000000000000001737177927613000000000000000000105851779050149", -- LUT(25) = log (0.9999999999999999999999996) = -1.7371779276130073106045160231020058517790501441178940472313536619042955E-25
		x"0000000000000000000000000173717792761300000000000000000017888143773428", -- LUT(26) = log (0.99999999999999999999999996) = -1.7371779276130073106045157104099788814377342353049807042811164431524514E-26
		x"0000000000000000000000000017371779276130000000000000000001761844036027", -- LUT(27) = log (0.999999999999999999999999996) = -1.7371779276130073106045156791407761844036026444236976250556047382880070E-27
		x"0000000000000000000000000001737177927613000000000000000000155914700186", -- LUT(28) = log (0.9999999999999999999999999996) = -1.7371779276130073106045156760138559147001894853355693996837486879716699E-28
		x"0000000000000000000000000000173717792761300000000000000000016388772985", -- LUT(29) = log (0.99999999999999999999999999996) = -1.7371779276130073106045156757011638877298481694267565779720700341417373E-29
		x"0000000000000000000000000000017371779276130000000000000000001946850324", -- LUT(30) = log (0.999999999999999999999999999996) = -1.7371779276130073106045156756698946850328140378358752958091572382707610E-30
		x"0000000000000000000000000000001737177927613000000000000000000167764763", -- LUT(31) = log (0.9999999999999999999999999999996) = -1.7371779276130073106045156756667677647631106246767871675929485093787836E-31
		x"0000000000000000000000000000000173717792761300000000000000000015507272", -- LUT(32) = log (0.99999999999999999999999999999996) = -1.7371779276130073106045156756664550727361402833608783547713284619965370E-32
		x"0000000000000000000000000000000017371779276130000000000000000001238031", -- LUT(33) = log (0.999999999999999999999999999999996) = -1.7371779276130073106045156756664238035334432492292874734891664655133819E-33
		x"0000000000000000000000000000000001737177927613000000000000000000120670", -- LUT(34) = log (0.9999999999999999999999999999999996) = -1.7371779276130073106045156756664206766131735458161283853609502659476171E-34
		x"0000000000000000000000000000000000173717792761300000000000000000012032", -- LUT(35) = log (0.99999999999999999999999999999999996) = -1.7371779276130073106045156756664203639211465754748124765481286459918661E-35
		x"0000000000000000000000000000000000017371779276130000000000000000001203"); -- LUT(36) = log (0.999999999999999999999999999999999996) = -1.7371779276130073106045156756664203639211465754748124765481286459918661E-36
	
signal lut_LogShP5: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"3010299956639800051200000000000130267681898814621085413104274611271087", -- LUT(1) = log (0.5) = -0.30102999566398119521373889472449302676818988146210854131042746112710819
		x"0222763947111520005120000000000017088170605440676109424036085924193578", -- LUT(2) = log (0.95) = -0.022276394711152233677405418967563708817060544067610942403608592419357348
		x"0021769192542745000000000000000001852733011099638352981197209562718919", -- LUT(3) = log (0.995) = -0.0021769192542745451137171103046901852733011099638352981197209562718910340
		x"0002172015458642500076800000000000167228838134068570615204766672430844", -- LUT(4) = log (0.9995) = -0.00021720154586425579969122400360587672288381340685706152047666724308432134
		x"0000217152669813610002560000000000016589513193002208080155018414844053", -- LUT(5) = log (0.99995) = -0.000021715266981361252472249012649395658951319300220808015501841484405957211
		x"0000021714778382153000000000000000001765705524336888830662761781040772", -- LUT(6) = log (0.999995) = -0.0000021714778382153786001749099590785765705524336888830662761781040778882661
		x"0000002171472952384500051200000000000161554391927873507132116189500642", -- LUT(7) = log (0.9999995) = -2.1714729523845424734224140533631615543919278735071321161895006417822643E-7
		x"0000000217147246380300007680000000000013387947451247399821039519863481", -- LUT(8) = log (0.99999995) = -2.1714724638030711857225321730389338794745124739982103951986348876620716E-8
		x"0000000021714724149449000768000000000001427855437372368866778314813782", -- LUT(9) = log (0.999999995) = -2.1714724149449401801418959207161427855437372368866778314813787638977192E-9
		x"0000000002171472410059100025600000000000150001130238267968999757062843", -- LUT(10) = log (0.9999999995) = -2.1714724100591272408156654133411500011302382679689997570628435304069588E-10
		x"0000000000217147240957050002560000000000014793413124046557253414145564", -- LUT(11) = log (0.99999999995) = -2.1714724095705459484953606333807479341312404655725341414556454303698637E-11
		x"0000000000021714724095216000000000000000001772263097741872398331067025", -- LUT(12) = log (0.999999999995) = -2.1714724095216878192794533380320772263097741872398331067028006293291233E-12
		x"0000000000002171472409516800000000000000000123449043417486138993950226", -- LUT(13) = log (0.9999999999995) = -2.1714724095168020063580238403236234490434174861389939502239156464987519E-13
		x"0000000000000217147240951630000000000000000014214385046674504612084487", -- LUT(14) = log (0.99999999999995) = -2.1714724095163134250658825028710421438504667450461208448295932178324262E-14
		x"0000000000000021714724095162000512000000000001666539961070472591713468", -- LUT(15) = log (0.999999999999995) = -2.1714724095162645669366683852489666539961070472591713462064028446304160E-15
		x"0000000000000002171472409516200076800000000000190931417260029770732189", -- LUT(16) = log (0.9999999999999995) = -2.1714724095162596811237469736479909314172600297707321817487912144107142E-16
		x"0000000000000000217147240951620007680000000000010567742344115714331780", -- LUT(17) = log (0.99999999999999995) = -2.1714724095162591925424548324895056774234411571433178555885208435762717E-17
		x"0000000000000000021714724095162000256000000000001732752066999281113899", -- LUT(18) = log (0.999999999999999995) = -2.1714724095162591436843256183736732752066999281113892459077825739501321E-18
		x"0000000000000000002171472409516200025600000000000190196216852211790448", -- LUT(19) = log (0.9999999999999999995) = -2.1714724095162591387985126969620901962168522117904441116960940687632083E-19
		x"0000000000000000000217147240951620002560000000000013188993018570422416", -- LUT(20) = log (0.99999999999999999995) = -2.1714724095162591383099314048209318899301857042241720151410161038963981E-20
		x"0000000000000000000021714724095162000256000000000001160593176422361087", -- LUT(21) = log (0.999999999999999999995) = -2.1714724095162591382610732756068160593176422361082030295937677432986701E-21
		x"0000000000000000000002171472409516200025600000000000104476256549121125", -- LUT(22) = log (0.9999999999999999999995) = -2.1714724095162591382561874626854044762565491211230127132800651001248192E-22
		x"0000000000000000000000217147240951620002560000000000016331795044142193", -- LUT(23) = log (0.99999999999999999999995) = -2.1714724095162591382556988813932633179504414219427577474711049973348204E-23
		x"0000000000000000000000021714724095162000256000000000001492021198306682", -- LUT(24) = log (0.999999999999999999999995) = -2.1714724095162591382556500232640492021198306681479148915484330886106929E-24
		x"0000000000000000000000002171472409516200025600000000000127790536769594", -- LUT(25) = log (0.9999999999999999999999995) = -2.1714724095162591382556451374511277905367695929296624323627481387537685E-25
		x"0000000000000000000000000217147240951620002560000000000013564937846341", -- LUT(26) = log (0.99999999999999999999999995) = -2.1714724095162591382556446488698356493784634854094495047082454661782309E-26
		x"0000000000000000000000000021714724095162000256000000000001064352626320", -- LUT(27) = log (0.999999999999999999999999995) = -2.1714724095162591382556446000117064352626328746574443351254358571447786E-27
		x"0000000000000000000000000002171472409516200025600000000000193513851040", -- LUT(28) = log (0.9999999999999999999999999995) = -2.1714724095162591382556445951258935138510498135822439793989813028236744E-28
		x"0000000000000000000000000000217147240951620002560000000000011222170980", -- LUT(29) = log (0.99999999999999999999999999995) = -2.1714724095162591382556445946373122217098915074747239454386541114573864E-29
		x"0000000000000000000000000000021714724095162000256000000000001540924950", -- LUT(30) = log (0.999999999999999999999999999995) = -2.1714724095162591382556445945884540924957756768639719420587445749614158E-30
		x"0000000000000000000000000000002171472409516200025600000000000168279573", -- LUT(31) = log (0.9999999999999999999999999999995) = -2.1714724095162591382556445945835682795743640938028967417209148531382254E-31
		x"0000000000000000000000000000000217147240951620002560000000000017969823", -- LUT(32) = log (0.99999999999999999999999999999995) = -2.1714724095162591382556445945830796982822229354967892216871334932741704E-32
		x"0000000000000000000000000000000021714724095162000256000000000001308403", -- LUT(33) = log (0.999999999999999999999999999999995) = -2.1714724095162591382556445945830308401530088196661784696837553734109475E-33
		x"0000000000000000000000000000000002171472409516200025600000000000125958", -- LUT(34) = log (0.9999999999999999999999999999999995) = -2.1714724095162591382556445945830259543400874080831173944834175615858571E-34
		x"0000000000000000000000000000000000217147240951620002560000000000012547", -- LUT(35) = log (0.99999999999999999999999999999999995) = -2.1714724095162591382556445945830254657587952669248112869633837804049603E-35
		x"0000000000000000000000000000000000021714724095162000256000000000001254"); -- LUT(36) = log (0.999999999999999999999999999999999995) = -2.1714724095162591382556445945830254657587952669248112869633837804049603E-36

signal lut_LogShP6: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"3979400086720300076800000000000139464636202370757829173791450777457830", -- LUT(1) = log (0.4) = -0.39794000867203760957252221055101394646362023707578291737914507774578362
		x"0268721464003010002560000000000013330720070201079436316522430875823190", -- LUT(2) = log (0.94) = -0.026872146400301340372041705826306333072007020107943631652243087582319967
		x"0026136156026866000768000000000001444778178206135340759092877140232678", -- LUT(3) = log (0.994) = -0.0026136156026866879812154116474416444778178206135340759092877140232674810
		x"0002606548934319700076800000000000110599250472668683015979854340416539", -- LUT(4) = log (0.9994) = -0.00026065489343197427769404564845954105992504726686830159798543404165379410
		x"0000260584506755330002560000000000014349920925528720185299613055230399", -- LUT(5) = log (0.99994) = -0.000026058450675533145391057860367025434992092552872018529961305523039353292
		x"0000026057747087514000512000000000001916302074430818495604938145289958", -- LUT(6) = log (0.999994) = -0.0000026057747087514545678487929202199916302074430818495604938145289954818797
		x"0000002605767673149800076800000000000158544986120740992357947451351187", -- LUT(7) = log (0.9999994) = -2.6057676731498910839277451065257585449861207409923579474513511893445724E-7
		x"0000000260576696959250002560000000000018578859593879205919041471441846", -- LUT(8) = log (0.99999994) = -2.6057669695925208354125129055348857885959387920591904147144184535039896E-8
		x"0000000026057668992368000512000000000001954372149294700936321658599335", -- LUT(9) = log (0.999999994) = -2.6057668992368116714345092489654954372149294700936321658599333896827449E-9
		x"0000000002605766892201200025600000000000115275929279074590199899280734", -- LUT(10) = log (0.9999999994) = -2.6057668922012410336453188303827152759292790745901998992807366490241337E-10
		x"0000000000260576689149760005120000000000017782374260248559113227717345", -- LUT(11) = log (0.99999999994) = -2.6057668914976839726524857627466778237426024855911322771734440950776161E-11
		x"0000000000026057668914273000512000000000001479891498839449144674755826", -- LUT(12) = log (0.999999999994) = -2.6057668914273282665810633156000479891498839449144674755821979390040453E-12
		x"0000000000002605766891420200076800000000000129496302459244919672064881", -- LUT(13) = log (0.9999999999994) = -2.6057668914202926959741996794814294963024592449196720648896199480039934E-13
		x"0000000000000260576689141950002560000000000012796667534089423707726462", -- LUT(14) = log (0.99999999999994) = -2.6057668914195891389135161019555279666753408942370772646936306998261860E-14
		x"0000000000000026057668914195000768000000000001974167839568060157741143", -- LUT(15) = log (0.999999999999994) = -2.6057668914195187832074477720637974167839568060157741146490903046626002E-15
		x"0000000000000002605766891419500025600000000000132957825406426167767754", -- LUT(16) = log (0.9999999999999994) = -2.6057668914195117476368409393532329578254064261677677515596067609547025E-16
		x"0000000000000000260576689141950002560000000000016259788985714322421403", -- LUT(17) = log (0.99999999999999994) = -2.6057668914195110440797802560849625978898571432242140092185365968106754E-17
		x"0000000000000000026057668914195000512000000000001634227559052723550222", -- LUT(18) = log (0.999999999999999994) = -2.6057668914195109737240741877581634227559052723550226095785631021103448E-18
		x"0000000000000000002605766891419500051200000000000183783851106115842222", -- LUT(19) = log (0.9999999999999999994) = -2.6057668914195109666885035809254837838511061158422298608661615431983970E-19
		x"0000000000000000000260576689141950005120000000000011582274671216049662", -- LUT(20) = log (0.99999999999999999994) = -2.6057668914195109659849465202422158227467121604966917246589429996681841E-20
		x"0000000000000000000026057668914195000512000000000001890266641336245655", -- LUT(21) = log (0.999999999999999999994) = -2.6057668914195109659145908141738890266641336245651953222996128670932280E-21
		x"0000000000000000000002605766891419500051200000000000156347056154379562", -- LUT(22) = log (0.9999999999999999999994) = -2.6057668914195109659075552435670563470561543795680762561761685225591675E-22
		x"0000000000000000000000260576689141950005120000000000017307909535924119", -- LUT(23) = log (0.99999999999999999999994) = -2.6057668914195109659068516865063730790953592411543246553049488495445015E-23
		x"0000000000000000000000026057668914195000512000000000001047522992797558", -- LUT(24) = log (0.999999999999999999999994) = -2.6057668914195109659067813308003047522992797551738090982752381297321738E-24
		x"0000000000000000000000002605766891419500051200000000000197919619671807", -- LUT(25) = log (0.9999999999999999999999994) = -2.6057668914195109659067742952296979196196718068543661386028411702257072E-25
		x"0000000000000000000000000260576689141950005120000000000013723635171105", -- LUT(26) = log (0.99999999999999999999999994) = -2.6057668914195109659067735916726372363517110120252079285959072153998080E-26
		x"0000000000000000000000000026057668914195000512000000000001311680249144", -- LUT(27) = log (0.999999999999999999999999994) = -2.6057668914195109659067735213169311680249149325423199684548168773284656E-27
		x"0000000000000000000000000002605766891419500051200000000000160561192233", -- LUT(28) = log (0.9999999999999999999999999994) = -2.6057668914195109659067735142813605611922353245940314510493038740954438E-28
		x"0000000000000000000000000000260576689141950005120000000000010350050892", -- LUT(29) = log (0.99999999999999999999999999994) = -2.6057668914195109659067735135778035005089673637992026020948385340778828E-29
		x"0000000000000000000000000000026057668914195000512000000000001477944401", -- LUT(30) = log (0.999999999999999999999999999994) = -2.6057668914195109659067735135074477944406405677197197172272528596791841E-30
		x"0000000000000000000000000000002605766891419500051200000000000112223831", -- LUT(31) = log (0.9999999999999999999999999999994) = -2.6057668914195109659067735135004122238338078881117714287407729008353448E-31
		x"0000000000000000000000000000000260576689141950005120000000000010866677", -- LUT(32) = log (0.99999999999999999999999999999994) = -2.6057668914195109659067735134997086667731246201509765998921276910369212E-32
		x"0000000000000000000000000000000026057668914195000512000000000001383116", -- LUT(33) = log (0.999999999999999999999999999999994) = -2.6057668914195109659067735134996383110670562933548971170072631979179384E-33
		x"0000000000000000000000000000000002605766891419500051200000000000131274", -- LUT(34) = log (0.9999999999999999999999999999999994) = -2.6057668914195109659067735134996312754964494606752891687187767488846487E-34
		x"0000000000000000000000000000000000260576689141950005120000000000013053", -- LUT(35) = log (0.99999999999999999999999999999999994) = -2.6057668914195109659067735134996305719393887774073283738899281039841058E-35
		x"0000000000000000000000000000000000026057668914195000512000000000001305"); -- LUT(36) = log (0.999999999999999999999999999999999994) = -2.6057668914195109659067735134996305719393887774073283738899281039841058E-36
signal lut_LogShP7: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"5228787452803300025600000000000146907998711358093041351701343596947709", -- LUT(1) = log (0.3) = -0.52287874528033756270497209674488469079987113580930413517013435969477085
		x"0315170514460640000000000000000019684961695775051194792317846396191807", -- LUT(2) = log (0.93) = -0.031517051446064883038267996626468968496169577505119479231784639619180240
		x"0030507515046188000768000000000001557171575861131595264405833674156596", -- LUT(3) = log (0.993) = -0.0030507515046188240968314894040280557171575861131595264405833674156592420
		x"0003041125891607600025600000000000188143439710191984843517576697050450", -- LUT(4) = log (0.9993) = -0.00030411258916076147349714559766534881434397101919848435175766970504586461
		x"0000304016778043650005120000000000013045937577925154454072651613680560", -- LUT(5) = log (0.99993) = -0.000030401677804365233665448449530405304593757792515445407265161368056137984
		x"0000030400720135872000000000000000001769224287622716499742625425239873", -- LUT(6) = log (0.999993) = -0.0000030400720135872240196786742857836769224287622716499742625425239873827181
		x"0000003040062437344700000000000000000193926217448196193093601935486192", -- LUT(7) = log (0.9999993) = -3.0400624373447400001432083043512939262174481961930936019354861980462508E-7
		x"0000000304006147972490000000000000000011099101214588912419389247093771", -- LUT(8) = log (0.99999993) = -3.0400614797249158252884373193994109910121458891241938924709377405625348E-8
		x"0000000030400613839629000256000000000001506065610661525363687271048736", -- LUT(9) = log (0.999999993) = -3.0400613839629776498419082348259506065610661525363687271048733186177025E-9
		x"0000000003040061374386700051200000000000104613262662879654630159923245", -- LUT(10) = log (0.9999999993) = -3.0400613743867842747174127680649046132626628796546301599232499232137729E-10
		x"0000000000304006137342910002560000000000015002568760221837833621827634", -- LUT(11) = log (0.99999999993) = -3.0400613734291649416291645637674500256876022183783362182763468288957927E-11
		x"0000000000030400613733334000000000000000001527670517934081016885070263", -- LUT(12) = log (0.999999999993) = -3.0400613733334030083645817565294527670517934081016885070260152974975160E-12
		x"0000000000003040061373323800000000000000000138484890732933630590756744", -- LUT(13) = log (0.9999999999993) = -3.0400613733238268150385658959373384848907329336305907567452767329815009E-13
		x"0000000000000304006137332280007680000000000014367907335352361149783783", -- LUT(14) = log (0.99999999999993) = -3.0400613733228691957059687340794436790733535236114978378553721261993612E-14
		x"0000000000000030400613733227000256000000000001673644835645504302240114", -- LUT(15) = log (0.999999999999993) = -3.0400613733227734337727090621356673644835645504302240110189865714625183E-15
		x"0000000000000003040061373322700051200000000000109864684273104491750633", -- LUT(16) = log (0.9999999999999993) = -3.0400613733227638575793830953837098646842731044917506375668957418195667E-16
		x"0000000000000000304006137332270007680000000000013831602094060237340122", -- LUT(17) = log (0.99999999999999993) = -3.0400613733227628999600504987129383160209406023734012880985116108349481E-17
		x"0000000000000000030400613733227000000000000000001054031677733183542831", -- LUT(18) = log (0.999999999999999993) = -3.0400613733227628041981172390459054031677733183542830344782389495763088E-18
		x"0000000000000000003040061373322700076800000000000102554302588249614069", -- LUT(19) = log (0.9999999999999999993) = -3.0400613733227627946219239130792025543025882496140663376309251397704477E-19
		x"0000000000000000000304006137332270007680000000000013227384027105933668", -- LUT(20) = log (0.99999999999999999993) = -3.0400613733227627936643045804825322738402710593366613871930423411519931E-20
		x"0000000000000000000030400613733227000768000000000001652458382813534747", -- LUT(21) = log (0.999999999999999999993) = -3.0400613733227627935685426472228652458382813534748870591096842485615679E-21
		x"0000000000000000000003040061373322700076800000000000198543038524803026", -- LUT(22) = log (0.9999999999999999999993) = -3.0400613733227627935589664538968985430385248030203692879707207028766874E-22
		x"0000000000000000000000304006137332270007680000000000010187275855357215", -- LUT(23) = log (0.99999999999999999999993) = -3.0400613733227627935580088345643018727585535721762341074735178389056424E-23
		x"0000000000000000000000030400613733227000768000000000001422057305564934", -- LUT(24) = log (0.999999999999999999999993) = -3.0400613733227627935579130726310422057305564933338337553899644871824741E-24
		x"0000000000000000000000003040061373322700076800000000000116239027756783", -- LUT(25) = log (0.9999999999999999999999993) = -3.0400613733227627935579034964377162390277567858920138518412708213566646E-25
		x"0000000000000000000000000304006137332270007680000000000018364235747682", -- LUT(26) = log (0.99999999999999999999999993) = -3.0400613733227627935579025388183836423574768151522560628029980714675484E-26
		x"0000000000000000000000000030400613733227000768000000000001503826904482", -- LUT(27) = log (0.999999999999999999999999993) = -3.0400613733227627935579024430564503826904488180783245259123367626455715E-27
		x"0000000000000000000000000003040061373322700076800000000000157056723742", -- LUT(28) = log (0.9999999999999999999999999993) = -3.0400613733227627935579024334802570567237460183709318146434022914250431E-28
		x"0000000000000000000000000000304006137332270007680000000000013772412701", -- LUT(29) = log (0.99999999999999999999999999993) = -3.0400613733227627935579024325226377241270757384001925479407101608996070E-29
		x"0000000000000000000000000000030400613733227000768000000000001757908672", -- LUT(30) = log (0.999999999999999999999999999993) = -3.0400613733227627935579024324268757908674087104031186213146829610130295E-30
		x"0000000000000000000000000000003040061373322700076800000000000199597543", -- LUT(31) = log (0.9999999999999999999999999999993) = -3.0400613733227627935579024324172995975414420076034112286525226611560315E-31
		x"0000000000000000000000000000000304006137332270007680000000000014197824", -- LUT(32) = log (0.99999999999999999999999999999993) = -3.0400613733227627935579024324163419782088453373234404893863110553716482E-32
		x"0000000000000000000000000000000030400613733227000768000000000001462165", -- LUT(33) = log (0.999999999999999999999999999999993) = -3.0400613733227627935579024324162462162755856702954434154596899390352231E-33
		x"0000000000000000000000000000000003040061373322700076800000000000136646", -- LUT(34) = log (0.9999999999999999999999999999999993) = -3.0400613733227627935579024324162366400822597035926437080670278278440007E-34
		x"0000000000000000000000000000000000304006137332270007680000000000013567", -- LUT(35) = log (0.99999999999999999999999999999999993) = -3.0400613733227627935579024324162356824629271069223637373277616167293027E-35
		x"0000000000000000000000000000000000030400613733227000768000000000001356"); -- LUT(36) = log (0.999999999999999999999999999999999993) = -3.0400613733227627935579024324162356824629271069223637373277616167293027E-36

signal lut_LogShP8: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"6989700043360100025600000000000169732318101185378914586895725388728910", -- LUT(1) = log (0.2) = -0.69897000433601880478626110527550697323181011853789145868957253887289181
		x"0362121726544440005120000000000013967661092027396867291035395911310940", -- LUT(2) = log (0.92) = -0.036212172654444730704745098299824396766109202739686729103539591131094985
		x"0034883278458213000512000000000001438553490343852726375095129742888688", -- LUT(3) = log (0.992) = -0.0034883278458213442646014262591191438553490343852726375095129742888684459
		x"0003475746339209000051200000000000127056576364768523547927965794579988", -- LUT(4) = log (0.9992) = -0.00034757463392090231671842480402357270565763647685235479279657945799850577
		x"0000347449483687260005120000000000014537727045641966189864783182628458", -- LUT(5) = log (0.99992) = -0.000034744948368726275656226672587143453772704564196618986478318262845072415
		x"0000034743697527235000512000000000001568810471722560238301477172320338", -- LUT(6) = log (0.999992) = -0.0000034743697527235555615660668462652568810471722560238301477172320332661655
		x"0000003474357244969000000000000000000190396094149326836960405653876420", -- LUT(7) = log (0.9999992) = -3.4743572449690979079753792188195903960941493268369604056538764250210910E-7
		x"0000000347435599420020002560000000000018414587067316633211918408767310", -- LUT(8) = log (0.99999992) = -3.4743559942002562422092187327698841458706731663321191840876731335218402E-8
		x"0000000034743558691234000000000000000001969646014145988067355439096579", -- LUT(9) = log (0.999999992) = -3.4743558691234381162326818590414969646014145988067355439096576403799324E-9
		x"0000000003474355856615700051200000000000120534499788101420359573246709", -- LUT(10) = log (0.9999999992) = -3.4743558566157569640406331160427205344997881014203595732467033467316929E-10
		x"0000000000347435585536490005120000000000016212781656633144106562916350", -- LUT(11) = log (0.99999999992) = -3.4743558553649888554254838953394621278165663314410656291635866875841251E-11
		x"0000000000034743558552399000256000000000001553834566426735076454984110", -- LUT(12) = log (0.999999999992) = -3.4743558552399120446300095294092553834566426735076454984115312696070841E-12
		x"0000000000003474355855227400051200000000000140052890212590088577374416", -- LUT(13) = log (0.9999999999992) = -3.4743558552274043635511224983772400528902125900885773744199587652772342E-13
		x"0000000000000347435585522610007680000000000014817742517193618440257715", -- LUT(14) = log (0.99999999999992) = -3.4743558552261535954432403993296481774251719361844025771343187651454959E-14
		x"0000000000000034743558552260000000000000000001450860587368010953080874", -- LUT(15) = log (0.999999999999992) = -3.4743558552260285186324522554654450860587368010953080873809676237745574E-15
		x"0000000000000003474355855226000000000000000000130337883498129796171343", -- LUT(16) = log (0.9999999999999992) = -3.4743558552260160109513734417394303378834981297961713471432633325343655E-16
		x"0000000000000000347435585522600005120000000000013291867558791524126212", -- LUT(17) = log (0.99999999999999992) = -3.4743558552260147601832655603734329186755879152412621599390238957935995E-17
		x"0000000000000000034743558552260000256000000000001992173108930299156741", -- LUT(18) = log (0.999999999999999992) = -3.4743558552260146351064547722368992173108930299156741928465527484080557E-18
		x"0000000000000000003474355855226000000000000000000146507579984502744012", -- LUT(19) = log (0.9999999999999999992) = -3.4743558552260146225987736934232465075799845027440185785603449216519194E-19
		x"0000000000000000000347435585522600000000000000000018124321094925964043", -- LUT(20) = log (0.99999999999999999992) = -3.4743558552260146213480055855418812432109492596404616531088612916164028E-20
		x"0000000000000000000034743558552260000000000000000001447168400862914264", -- LUT(21) = log (0.999999999999999999992) = -3.4743558552260146212229287747537447168400862914262420465276372068990124E-21
		x"0000000000000000000003474355855226000000000000000000131064203660400165", -- LUT(22) = log (0.9999999999999999999992) = -3.4743558552260146212104210936749310642036604001657814467287581941168948E-22
		x"0000000000000000000000347435585522600000000000000000014969894002441507", -- LUT(23) = log (0.99999999999999999999992) = -3.4743558552260146212091703255670496989400244150953450003574623309484860E-23
		x"0000000000000000000000034743558552260000000000000000001615624136608827", -- LUT(24) = log (0.999999999999999999999992) = -3.4743558552260146212090452487562615624136608826288574518564186646168960E-24
		x"0000000000000000000000003474355855226000000000000000000182748761024537", -- LUT(25) = log (0.9999999999999999999999992) = -3.4743558552260146212090327410751827487610245300426142579676751571831937E-25
		x"0000000000000000000000000347435585522600000000000000000017486739576089", -- LUT(26) = log (0.99999999999999999999999992) = -3.4743558552260146212090314903070748673957608947905939941884144150318176E-26
		x"0000000000000000000000000034743558552260000000000000000001640792592348", -- LUT(27) = log (0.999999999999999999999999992) = -3.4743558552260146212090313652302640792592345312654580083665844769026000E-27
		x"0000000000000000000000000003474355855226000000000000000000183000445587", -- LUT(28) = log (0.9999999999999999999999999992) = -3.4743558552260146212090313527225830004455818949129450701899624444505374E-28
		x"0000000000000000000000000000347435585522600000000000000000011489256426", -- LUT(29) = log (0.99999999999999999999999999992) = -3.4743558552260146212090313514718148925642166312776937829763558508189397E-29
		x"0000000000000000000000000000034743558552260000000000000000001380817765", -- LUT(30) = log (0.999999999999999999999999999992) = -3.4743558552260146212090313513467380817760801049141686543210357475519161E-30
		x"0000000000000000000000000000003474355855226000000000000000000130400694", -- LUT(31) = log (0.9999999999999999999999999999992) = -3.4743558552260146212090313513342304006972664522778161414561641427861750E-31
		x"0000000000000000000000000000000347435585522600000000000000000017963251", -- LUT(32) = log (0.99999999999999999999999999999992) = -3.4743558552260146212090313513329796325893850870141808901696835863652106E-32
		x"0000000000000000000000000000000034743558552260000000000000000001545552", -- LUT(33) = log (0.999999999999999999999999999999992) = -3.4743558552260146212090313513328545557785969504878173650410355967636702E-33
		x"0000000000000000000000000000000003474355855226000000000000000000142041", -- LUT(34) = log (0.9999999999999999999999999999999992) = -3.4743558552260146212090313513328420480975181368351810125281707984639217E-34
		x"0000000000000000000000000000000000347435585522600000000000000000014071", -- LUT(35) = log (0.99999999999999999999999999999999992) = -3.4743558552260146212090313513328407973294102554699173772768843186405509E-35
		x"0000000000000000000000000000000000034743558552260000000000000000001407"); -- LUT(36) = log (0.999999999999999999999999999999999992) = -3.4743558552260146212090313513328407973294102554699173772768843186405509E-36

signal lut_LogShP9: mlut_LogShP := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2787536009528200000000000000000193179511293373944975989068188687077500", -- LUT(1) = log (0.1) = -1
		x"0409586076789060000000000000000013756866984152889663216951740712841936", -- LUT(2) = log (0.91) = -0.040958607678906400081278583465035375686698415288966321695174071284193468
		x"0039263455147246000256000000000001358674873367718791812151581960013847", -- LUT(3) = log (0.991) = -0.0039263455147246716355656211845791358674873367718791812151581960013842878
		x"0003910410285829400025600000000000161836349183851024605284713938485536", -- LUT(4) = log (0.9991) = -0.00039104102858294304456699375418312618363491838510246052847139384855318914
		x"0000390882623694850007680000000000012710397251821395083231460133433506", -- LUT(5) = log (0.99991) = -0.000039088262369485055789164769170025271039725182139508323146013343350606835
		x"0000039086679261613000000000000000001565591370816649292686345345616717", -- LUT(6) = log (0.999991) = -0.0000039086679261613178020183232463383565591370816649292686345345616713899101
		x"0000003908652096022900076800000000000150314699905425992182583130854206", -- LUT(7) = log (0.9999991) = -3.9086520960229734933334391960980503146999054259921825831308542007082972E-7
		x"0000000390865051301850005120000000000010094668817457954956510172756873", -- LUT(8) = log (0.99999991) = -3.9086505130185421730337730695513009466881745795495651017275687948069176E-8
		x"0000000039086503547181000512000000000001901467362273346613458778509122", -- LUT(9) = log (0.999999991) = -3.9086503547181930714754191049618901467362273346613458778509120410855037E-9
		x"0000000003908650338888100000000000000000171327908768816420193694408031", -- LUT(10) = log (0.9999999991) = -3.9086503388881591016236657639737713279087688164201936944080321320264795E-10
		x"0000000000390865033730510000000000000000011432374671364141193580702211", -- LUT(11) = log (0.99999999991) = -3.9086503373051557140415306163591143237467136414119358070221473420323320E-11
		x"0000000000039086503371468000512000000000001196644113387293309601859832", -- LUT(12) = log (0.999999999991) = -3.9086503371468553753773475028284196644113387293309601859838297523417705E-12
		x"0000000000003908650337131000025600000000000123838385478019001886073658", -- LUT(13) = log (0.9999999999991) = -3.9086503371310253415118694954870238383854780190018860736559415697364733E-13
		x"0000000000000390865033712940002560000000000010035811146604073770291559", -- LUT(14) = log (0.99999999999991) = -3.9086503371294423381253310977930003581114660407377029155905525212292394E-14
		x"0000000000000039086503371292000256000000000001991704732800812095802879", -- LUT(15) = log (0.999999999999991) = -3.9086503371292840377866773520539991704732800812095802872194933677228383E-15
		x"0000000000000003908650337129200000000000000000103063312719567137126159", -- LUT(16) = log (0.9999999999999991) = -3.9086503371292682077528119784204030633127195671371261545527342268902114E-16
		x"0000000000000000390865033712920000000000000000014649271269546247818161", -- LUT(17) = log (0.99999999999999991) = -3.9086503371292666247494254410664464927126954624781816982175428813428349E-17
		x"0000000000000000039086503371292000512000000000001448660538533708456991", -- LUT(18) = log (0.999999999999999991) = -3.9086503371292664664490867873311448660538533708456997595290140220851282E-18
		x"0000000000000000003908650337129200025600000000000115643691980764870152", -- LUT(19) = log (0.9999999999999999991) = -3.9086503371292664506190529219576156436919807648701516202269867189067906E-19
		x"0000000000000000000390865033712920002560000000000016273085883362030440", -- LUT(20) = log (0.99999999999999999991) = -3.9086503371292664490360495354202627308588336203044731727719496200968821E-20
		x"0000000000000000000039086503371292000256000000000001274396695493070080", -- LUT(21) = log (0.999999999999999999991) = -3.9086503371292664488777491967665274396695493070082240910571270639066510E-21
		x"0000000000000000000003908650337129200025600000000000153910551561179690", -- LUT(22) = log (0.9999999999999999999991) = -3.9086503371292664488619191629011539105515611796902023705153175493219112E-22
		x"0000000000000000000000390865033712920002560000000000011655763977176994", -- LUT(23) = log (0.99999999999999999999991) = -3.9086503371292664488603361595146165576397717699985162303374326912032774E-23
		x"0000000000000000000000039086503371292000256000000000001628223485929236", -- LUT(24) = log (0.999999999999999999999991) = -3.9086503371292664488601778591759628223485929230597487766384071656907419E-24
		x"0000000000000000000000003908650337129200025600000000000197448819475037", -- LUT(25) = log (0.9999999999999999999999991) = -3.9086503371292664488601620291420974488194750393061760428716922427418476E-25
		x"0000000000000000000000000390865033712920002560000000000011091146656328", -- LUT(26) = log (0.99999999999999999999999991) = -3.9086503371292664488601604461387109114665632509402218096110526267429811E-26
		x"0000000000000000000000000039086503371292000256000000000001722577312721", -- LUT(27) = log (0.999999999999999999999999991) = -3.9086503371292664488601602878383722577312720721037204166861489839060547E-27
		x"0000000000000000000000000003908650337129200025600000000000138392357741", -- LUT(28) = log (0.9999999999999999999999999991) = -3.9086503371292664488601602720083383923577429542200712176976702228099917E-28
		x"0000000000000000000000000000390865033712920002560000000000013500582036", -- LUT(29) = log (0.99999999999999999999999999991) = -3.9086503371292664488601602704253350058203900424317063072018624627322616E-29
		x"0000000000000000000000000000039086503371292000256000000000001346671667", -- LUT(30) = log (0.999999999999999999999999999991) = -3.9086503371292664488601602702670346671666547512528698162463120878848074E-30
		x"0000000000000000000000000000003908650337129200025600000000000104633307", -- LUT(31) = log (0.9999999999999999999999999999991) = -3.9086503371292664488601602702512046333012812221349861671516973544116652E-31
		x"0000000000000000000000000000000390865033712920002560000000000012162999", -- LUT(32) = log (0.99999999999999999999999999999991) = -3.9086503371292664488601602702496216299147438692231978022422452841044670E-32
		x"0000000000000000000000000000000039086503371292000256000000000001633298", -- LUT(33) = log (0.999999999999999999999999999999991) = -3.9086503371292664488601602702494633295760901339320189657513001711041483E-33
		x"0000000000000000000000000000000003908650337129200025600000000000147490", -- LUT(34) = log (0.9999999999999999999999999999999991) = -3.9086503371292664488601602702494474995422247604029010821022056607444205E-34
		x"0000000000000000000000000000000000390865033712920002560000000000014591", -- LUT(35) = log (0.99999999999999999999999999999999991) = -3.9086503371292664488601602702494459165388382230499892937372962097178507E-35
		x"0000000000000000000000000000000000039086503371292000256000000000001459"); -- LUT(36) = log (0.999999999999999999999999999999999991) = -3.9086503371292664488601602702494459165388382230499892937372962097178507E-36


-- ====== FIN declaraci�n
-- declaracion de meomria de log para la parte de x>1

-- ====== Comienzo declaraci�n
-- declaracion de meomria de log para la parte de x<1

type mlut_LogShN is array (0 to P+2) of std_logic_vector (8*P+7 downto 0);

signal lut_LogShN9: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"0413926851582250005120000000000012417067021904664530945965390186797530", -- LUT(1) = log (1.1) = 0.041392685158225040750199971243024241706702190466453094596539018679753032
		x"0043213737826425000512000000000001132192893552064525914058186369484480", -- LUT(2) = log (1.01) = 0.0043213737826425742751881782229379132192893552064525914058186369484480104
		x"0004340774793186400076800000000000160200037751774867729013649473955591", -- LUT(3) = log (1.001) = 0.00043407747931864066892138777798886602000377517748677290136494739555956377
		x"0000434272768626690002560000000000011310979627758925307732464042115841", -- LUT(4) = log (1.0001) = 0.000043427276862669637313527585098268131097962775892530773246404211584759011
		x"0000043429231044531000512000000000001839724439448249094541443880968620", -- LUT(5) = log (1.00001) = 0.0000043429231044531868554934716343971839724439448249094541443880968627435425
		x"0000004342942647561500000000000000000170416841361667145121612010092062", -- LUT(6) = log (1.000001) = 4.3429426475615564074394264367770704168413616671451216120100920600646163E-7
		x"0000000434294460188520000000000000000014716184534126294027719584836885", -- LUT(7) = log (1.0000001) = 4.3429446018852918013670197358779471618453412629402771958483688371187471E-8
		x"0000000043429447973177000256000000000001513552500188036530684122042806", -- LUT(8) = log (1.00000001) = 4.3429447973177943261135240219573513552500188036530684122042800710352334E-9
		x"0000000004342944816861000051200000000000109449975167103574888128566606", -- LUT(9) = log (1.000000001) = 4.3429448168610458684426783228355094499751671035748881285666077943342844E-10
		x"0000000000434294481881530002560000000000010902153603387684726625081276", -- LUT(10) = log (1.0000000001) = 4.3429448188153710355741397580695090215360338768472662508127253947631500E-11
		x"0000000000043429448190108000512000000000001943752044854307845718560527", -- LUT(11) = log (1.00000000001) = 4.3429448190108035524162713626107943752044854307845718560521428168814761E-12
		x"0000000000004342944819030300000000000000000168188103076331630995751301", -- LUT(12) = log (1.000000000001) = 4.3429448190303468041017743776760681881030763316309957513017772960244133E-13
		x"0000000000000434294481903230002560000000000010798859182027432839105041", -- LUT(13) = log (1.0000000000001) = 4.3429448190323011292703375777287079885918202743283910504849072998679919E-14
		x"0000000000000043429448190324000512000000000001330937991070845967224892", -- LUT(14) = log (1.00000000000001) = 4.3429448190324965617871940267194330937991070845967224894788994375775741E-15
		x"0000000000000004342944819032500000000000000000160215572386313351021740", -- LUT(15) = log (1.000000000000001) = 4.3429448190325161050388796729083602155723863133510217474644354630612721E-16
		x"0000000000000000434294481903250005120000000000015147386224070812729389", -- LUT(16) = log (1.0000000000000001) = 4.3429448190325180593640482375401514738622407081272938153719073538458377E-17
		x"0000000000000000043429448190325000512000000000001595851523514132903538", -- LUT(17) = log (1.00000000000000001) = 4.3429448190325182547965650940034595851523514132903530110647890888807852E-18
		x"0000000000000000004342944819032500051200000000000191686135973736464473", -- LUT(18) = log (1.000000000000000001) = 4.3429448190325182743398167796497916861359737364644796740905796609375344E-19
		x"0000000000000000000434294481903250005120000000000012490913288208130842", -- LUT(19) = log (1.0000000000000000001) = 4.3429448190325182762941419482144249091328820813084715142512912231826086E-20
		x"0000000000000000000043429448190325000512000000000001882315615583769180", -- LUT(20) = log (1.00000000000000000001) = 4.3429448190325182764895744650708882315615583769181364909723672719385639E-21
		x"0000000000000000000004342944819032500051200000000000134563805715861092", -- LUT(21) = log (1.000000000000000000001) = 4.3429448190325182765091177167565345638057158610903556465724913493069550E-22
		x"0000000000000000000000434294481903250005120000000000019919703014450801", -- LUT(22) = log (1.0000000000000000000001) = 4.3429448190325182765110720419250991970301445080536900887117848881922896E-23
		x"0000000000000000000000043429448190325000512000000000001556603525875011", -- LUT(23) = log (1.00000000000000000000001) = 4.3429448190325182765112674744419556603525875017354846581915070543587315E-24
		x"0000000000000000000000004342944819032500051200000000000141306684831808", -- LUT(24) = log (1.000000000000000000000001) = 4.3429448190325182765112870176936413066848318023935187263921371990991212E-25
		x"0000000000000000000000000434294481903250005120000000000010987131805629", -- LUT(25) = log (1.0000000000000000000000001) = 4.3429448190325182765112889720188098713180562324722206793247267928543986E-26
		x"0000000000000000000000000043429448190325000512000000000001267277813780", -- LUT(26) = log (1.00000000000000000000000001) = 4.3429448190325182765112891674513267277813786754802198600791110180227388E-27
		x"0000000000000000000000000004342944819032500051200000000000178413427719", -- LUT(27) = log (1.000000000000000000000000001) = 4.3429448190325182765112891869945784134277109197810210680091606931975009E-28
		x"0000000000000000000000000000434294481903250005120000000000010358199230", -- LUT(28) = log (1.0000000000000000000000000001) = 4.3429448190325182765112891889489035819923441442111012017007117732415564E-29
		x"0000000000000000000000000000043429448190325000512000000000001360988481", -- LUT(29) = log (1.00000000000000000000000000001) = 4.3429448190325182765112891891443360988488074666541092151988523423712277E-30
		x"0000000000000000000000000000004342944819032500051200000000000179350532", -- LUT(30) = log (1.000000000000000000000000000001) = 4.3429448190325182765112891891638793505344537988984100165499562538954475E-31
		x"0000000000000000000000000000000434294481903250005120000000000013367572", -- LUT(31) = log (1.0000000000000000000000000000001) = 4.3429448190325182765112891891658336757030184321228400966850795435939820E-32
		x"0000000000000000000000000000000043429448190325000512000000000001291083", -- LUT(32) = log (1.00000000000000000000000000000001) = 4.3429448190325182765112891891660291082198748954452831046985920015492966E-33
		x"0000000000000000000000000000000004342944819032500051200000000000148654", -- LUT(33) = log (1.000000000000000000000000000000001) = 4.3429448190325182765112891891660486514715605417775274054999432486346827E-34
		x"0000000000000000000000000000000000434294481903250005120000000000015065", -- LUT(34) = log (1.0000000000000000000000000000000001) = 4.3429448190325182765112891891660506057967291064107518355800783733561198E-35
		x"0000000000000000000000000000000000043429448190325000512000000000001506", -- LUT(35) = log (1.00000000000000000000000000000000001) = 4.3429448190325182765112891891660508012292459628740742785880918858283925E-36
		x"0000000000000000000000000000000000004342944819032500051200000000000150");-- LUT(36) = log (1.000000000000000000000000000000000001) = 4.3429448190325182765112891891660508012292459628740742785880918858283925E-37


signal lut_LogShN8: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"0791812460476240005120000000000013627365086271149129474507205625594450", -- LUT(1) = log (1.2) = 0.079181246047624827722505692704101362736508627114912947450720562559445531
		x"0086001717619175000256000000000001659758861240778508035206615837770319", -- LUT(2) = log (1.02) = 0.0086001717619175610489366923079453659758861240778508035206615837770314043
		x"0008677215312269100025600000000000104296571469840626350472566290986008", -- LUT(3) = log (1.002) = 0.00086772153122691249284270790007587042965714698406263504725662909860080774
		x"0000868502116489570007680000000000016291373319656945431149891112722667", -- LUT(4) = log (1.0002) = 0.000086850211648957228899798162210906629137331965694543114989111272266502517
		x"0000086858027803267000256000000000001427235713814461666611150027033256", -- LUT(5) = log (1.00002) = 0.0000086858027803267571495643873989012427235713814461666611150027033250175526
		x"0000008685880952186900051200000000000197455039912229762838045828539065", -- LUT(6) = log (1.000002) = 8.6858809521869796567983605898281974550399122297628380458285390641260595E-7
		x"0000000868588876947610005120000000000015826155021854587743163487365994", -- LUT(7) = log (1.0000002) = 8.6858887694761885583633921667316582615502185458774316348736599224486314E-8
		x"0000000086858895512061000256000000000001600839680536630928688321540233", -- LUT(8) = log (1.00000002) = 8.6858895512061413304908138849988600839680536630928688321540235051613215E-9
		x"0000000008685889629379100025600000000000159423250716664066408956808032", -- LUT(9) = log (1.000000002) = 8.6858896293791469265387279920244594232507166640664089568080317123699482E-10
		x"0000000000868588963719640007680000000000013918282168040810663774011991", -- LUT(10) = log (1.0000000002) = 8.6858896371964475893318865848533391828216804081066377401199340329905979E-11
		x"0000000000086858896379781000512000000000001671618657462579402585696390", -- LUT(11) = log (1.00000000002) = 8.6858896379781776566430861314202671618657462579402585696397326344071560E-12
		x"0000000000008685889638056300051200000000000163136853232768429669565772", -- LUT(12) = log (1.000000000002) = 8.6858896380563506633845249229652631368532327684296695657718018848092247E-13
		x"0000000000000868588963806410005120000000000016122889988916693366027903", -- LUT(13) = log (1.0000000000002) = 8.6858896380641679640587719904886612288998891669336602790841292989493843E-14
		x"0000000000000086858896380649000768000000000001900385128109636806067634", -- LUT(14) = log (1.00000000000002) = 8.6858896380649496941261977291246900385128109636806067635370375727171153E-15
		x"0000000000000008685889638065000051200000000000129809493648482003936265", -- LUT(15) = log (1.000000000000002) = 8.6858896380650278671329403133071298094936484820039362627233570809821730E-16
		x"0000000000000000868588963806500007680000000000016215549194314999983526", -- LUT(16) = log (1.0000000000000002) = 8.6858896380650356844336145718285621554919431499998352552639784136795455E-17
		x"0000000000000000086858896380650000512000000000001372737807747414238377", -- LUT(17) = log (1.00000000000000002) = 8.6858896380650364661636819976817372737807747414238378946408488167913711E-18
		x"0000000000000000008685889638065000025600000000000165104446547921827948", -- LUT(18) = log (1.000000000000000002) = 8.6858896380650365443366887402670651044465479218279450630594607755566908E-19
		x"0000000000000000000868588963806500005120000000000019799070149414008099", -- LUT(19) = log (1.0000000000000000002) = 8.6858896380650365521539894145255979907014941400809883117232109174782578E-20
		x"0000000000000000000086858896380650000512000000000001512803588724509082", -- LUT(20) = log (1.00000000000000000002) = 8.6858896380650365529357194819514512803588724509084189773705819008277278E-21
		x"0000000000000000000008685889638065000051200000000000136609334929118883", -- LUT(21) = log (1.000000000000000000002) = 8.6858896380650365530138924886940366093349291188811833073585917359339448E-22
		x"0000000000000000000000868588963806500005120000000000019514223263797405", -- LUT(22) = log (1.0000000000000000000002) = 8.6858896380650365530217097893682951422326379740473599529916409095893589E-23
		x"0000000000000000000000086858896380650000512000000000001209955224098913", -- LUT(23) = log (1.00000000000000000000002) = 8.6858896380650365530224915194357209955224098914476666196812883243191253E-24
		x"0000000000000000000000008685889638065000051200000000000163580851387094", -- LUT(24) = log (1.000000000000000000000002) = 8.6858896380650365530225696924424635808513870935065341763715164907812070E-25
		x"0000000000000000000000000868588963806500005120000000000013783938428484", -- LUT(25) = log (1.0000000000000000000000002) = 8.6858896380650365530225775097431378393842848138156093009407519416773217E-26
		x"0000000000000000000000000086858896380650000512000000000001052652375744", -- LUT(26) = log (1.00000000000000000000000002) = 8.6858896380650365530225782914732052652375745858475486970866776131094322E-27
		x"0000000000000000000000000008685889638065000051200000000000112007822900", -- LUT(27) = log (1.000000000000000000000000002) = 8.6858896380650365530225783696462120078229035630507529555381602015160683E-28
		x"0000000000000000000000000000868588963806500005120000000000011268208140", -- LUT(28) = log (1.0000000000000000000000000002) = 8.6858896380650365530225783774635126820814364607710734845716773605693661E-29
		x"0000000000000000000000000000086858896380650000512000000000001427495070", -- LUT(29) = log (1.00000000000000000000000000002) = 8.6858896380650365530225783782452427495072897505431055385069127654768223E-30
		x"0000000000000000000000000000008685889638065000051200000000000115756240", -- LUT(30) = log (1.000000000000000000000000000002) = 8.6858896380650365530225783783234157562498750795203087439107551428575891E-31
		x"0000000000000000000000000000000868588963806500005120000000000013305698", -- LUT(31) = log (1.0000000000000000000000000000002) = 8.6858896380650365530225783783312330569241336124180290644512425689645660E-32
		x"0000000000000000000000000000000086858896380650000512000000000001147868", -- LUT(32) = log (1.00000000000000000000000000000002) = 8.6858896380650365530225783783320147869915594657078010965052923434589527E-33
		x"0000000000000000000000000000000008685889638065000051200000000000192959", -- LUT(33) = log (1.000000000000000000000000000000002) = 8.6858896380650365530225783783320929599983020510367782997106973312272283E-34
		x"0000000000000000000000000000000000868588963806500005120000000000010075", -- LUT(34) = log (1.0000000000000000000000000000000002) = 8.6858896380650365530225783783321007772989763095696760200312378301072442E-35
		x"0000000000000000000000000000000000086858896380650000512000000000001014", -- LUT(35) = log (1.00000000000000000000000000000000002) = 8.6858896380650365530225783783321015590290437354229657920632918799962777E-36
		x"0000000000000000000000000000000000008685889638065000051200000000000101"); -- LUT(36) = log (1.000000000000000000000000000000000002) = 8.6858896380650365530225783783321015590290437354229657920632918799962777E-37


signal lut_LogShN7: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"1139433523068300076800000000000184308297291883870682718011909749975530", -- LUT(1) = log (1.3) = 0.11394335230683676920650515794232843082972918838706827180119097499755309
		x"0128372247051720000000000000000014243905234969760305647528079332618920", -- LUT(2) = log (1.03) = 0.012837224705172205171071194580239424390523496976030564752807933261892818
		x"0013009330204181000000000000000001689343118533558116129076540476281440", -- LUT(3) = log (1.003) = 0.0013009330204181188008262788634812689343118533558116129076540476281448091
		x"0001302688052270600025600000000000181134370779944226787491282936416642", -- LUT(4) = log (1.0003) = 0.00013026880522706100378087172925158811343707799442267874912829364166466392
		x"0000130286390284890005120000000000017779794526944078367167882625656712", -- LUT(5) = log (1.00003) = 0.000013028639028489260760818724016476777979452694407836716788262565671367474
		x"0000013028814913884000512000000000001446266684366636420812809974702753", -- LUT(6) = log (1.000003) = 0.0000013028814913884955598628494412367446266684366636420812809974702754565810
		x"0000001302883250277200000000000000000120140885815174684151057156755064", -- LUT(7) = log (1.0000003) = 1.3028832502772777129846411452584201408858151746841510571567550647001717E-7
		x"0000000130288342616650007680000000000011130791540770631590038082997395", -- LUT(8) = log (1.00000003) = 1.3028834261665041881720794309126113079154077063159003808299739003801761E-8
		x"0000000013028834437554000000000000000001383231844906751315577131009546", -- LUT(9) = log (1.000000003) = 1.3028834437554303182974038606545383231844906751315577131009545416576293E-9
		x"0000000001302883445514300051200000000000105434602890154752602278617157", -- LUT(10) = log (1.0000000003) = 1.3028834455143229661360099376693054346028901547526022786171535939318215E-10
		x"0000000000130288344569020002560000000000011857771357147495238504199938", -- LUT(11) = log (1.00000000003) = 1.3028834456902122312681312895392185777135714749523850419993635335345813E-11
		x"0000000000013028834457078000512000000000001222872200518961812023631488", -- LUT(12) = log (1.000000000003) = 1.3028834457078011577848260321757222872200518961812023631480701635061720E-12
		x"0000000000001302883445709500025600000000000175610153548570467031183341", -- LUT(13) = log (1.0000000000003) = 1.3028834457095600504365303325138756101535485704670311833464537947067263E-13
		x"0000000000000130288344570970002560000000000013597979475762060505393682", -- LUT(14) = log (1.00000000000003) = 1.3028834457097359397017011108084359797947576206050539368646019414114432E-14
		x"0000000000000013028834457097000256000000000001994671401851503425262753", -- LUT(15) = log (1.000000000000003) = 1.3028834457097535286282181921204994671401851503425262752862562755151559E-15
		x"0000000000000001302883445709700076800000000000131890378548797594406801", -- LUT(16) = log (1.0000000000000003) = 1.3028834457097552875208699002865318903785487975944068042088703849057815E-16
		x"0000000000000000130288344570970005120000000000018339344742337909040702", -- LUT(17) = log (1.00000000000000003) = 1.3028834457097554634101350711034833934474233790904070866482645724278737E-17
		x"0000000000000000013028834457097000768000000000001820263617612194155431", -- LUT(18) = log (1.000000000000000003) = 1.3028834457097554809990615881851820263617612194155432680842718350896907E-18
		x"0000000000000000001302883445709700076800000000000151924479269507269821", -- LUT(19) = log (1.0000000000000000003) = 1.3028834457097554827579542398933519244792695072698200757906898363298976E-19
		x"0000000000000000000130288344570970007680000000000016891463928108109342", -- LUT(20) = log (1.00000000000000000003) = 1.3028834457097554829338435050641689146392810810934653962849907058001954E-20
		x"0000000000000000000013028834457097000768000000000001506136587648459265", -- LUT(21) = log (1.000000000000000000003) = 1.3028834457097554829514324315812506136587648459262121047394854143372844E-21
		x"0000000000000000000001302883445709700076800000000000158783560748048486", -- LUT(22) = log (1.0000000000000000000003) = 1.3028834457097554829531913242329587835607480484839905973489933594377905E-22
		x"0000000000000000000000130288344570970007680000000000012960055094671707", -- LUT(23) = log (1.00000000000000000000003) = 1.3028834457097554829533672134981296005509467170005134848275847465183400E-23
		x"0000000000000000000000013028834457097000768000000000001466822499665875", -- LUT(24) = log (1.000000000000000000000003) = 1.3028834457097554829533848024246466822499665873347732239576202911599280E-24
		x"0000000000000000000000001302883445709700076800000000000198390419868574", -- LUT(25) = log (1.0000000000000000000000003) = 1.3028834457097554829533865613172983904198685744030252723744456096834299E-25
		x"0000000000000000000000000130288344570970007680000000000016356123685872", -- LUT(26) = log (1.00000000000000000000000003) = 1.3028834457097554829533867372065635612368587731101987379611663591763736E-26
		x"0000000000000000000000000013028834457097000768000000000001900783185571", -- LUT(27) = log (1.000000000000000000000000003) = 1.3028834457097554829533867547954900783185577929809195671272888163020739E-27
		x"0000000000000000000000000001302883445709700076800000000000182730026729", -- LUT(28) = log (1.0000000000000000000000000003) = 1.3028834457097554829533867565543827300267276949679916848699755658364080E-28
		x"0000000000000000000000000000130288344570970007680000000000017199519758", -- LUT(29) = log (1.00000000000000000000000000003) = 1.3028834457097554829533867567302719951975446851666988969925049858280590E-29
		x"0000000000000000000000000000013028834457097000768000000000001609217144", -- LUT(30) = log (1.000000000000000000000000000003) = 1.3028834457097554829533867567478609217146263841865696182082405352776063E-30
		x"0000000000000000000000000000001302883445709700076800000000000119814363", -- LUT(31) = log (1.0000000000000000000000000000003) = 1.3028834457097554829533867567496198143663345540885566903298489162970648E-31
		x"0000000000000000000000000000000130288344570970007680000000000019570363", -- LUT(32) = log (1.00000000000000000000000000000003) = 1.3028834457097554829533867567497957036315053710787553975420101026597557E-32
		x"0000000000000000000000000000000013028834457097000768000000000001132923", -- LUT(33) = log (1.000000000000000000000000000000003) = 1.3028834457097554829533867567498132925580224527777752682632262247786323E-33
		x"0000000000000000000000000000000001302883445709700076800000000000115055", -- LUT(34) = log (1.0000000000000000000000000000000003) = 1.3028834457097554829533867567498150514506741609476772553353478370253460E-34
		x"0000000000000000000000000000000000130288344570970007680000000000011525", -- LUT(35) = log (1.00000000000000000000000000000000003) = 1.3028834457097554829533867567498152273399393317646674540425599982503656E-35
		x"0000000000000000000000000000000000013028834457097000768000000000001152"); -- LUT(36) = log (1.000000000000000000000000000000000003) = 1.3028834457097554829533867567498152273399393317646674540425599982503656E-36

signal lut_LogShN6: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"1461280356782300051200000000000192202517622777860739478140624148453610", -- LUT(1) = log (1.4) = 0.14612803567823802592595515331712922025176227778607394781406241484536163
		x"0170333392987800007680000000000015111342988327733938957324733583788779", -- LUT(2) = log (1.04) = 0.017033339298780354847721842115807511134298832773393895732473358378877659
		x"0017337128090005000512000000000001353938464483173693912766526348677875", -- LUT(3) = log (1.004) = 0.0017337128090005297680271061558901353938464483173693912766526348677872180
		x"0001736830584649100025600000000000123302721538713083836985606118111005", -- LUT(4) = log (1.0004) = 0.00017368305846491882263815317448820233027215387130838369856061181110027797
		x"0000173714318498090005120000000000013584970364956774925459314230068555", -- LUT(5) = log (1.00004) = 0.000017371431849809221512278044616760358497036495677492545931423006855061444
		x"0000017371744532664000000000000000001925464236143372274419302357944895", -- LUT(6) = log (1.000004) = 0.0000017371744532664170057424059403635925464236143372274419302357944893341770
		x"0000001737177580177500025600000000000157344355836280300086931476653715", -- LUT(7) = log (1.0000004) = 1.7371775801775144374647314105390573443558362803000869314766537195320619E-7
		x"0000000173717789286940007680000000000018676520986214696453543976270605", -- LUT(8) = log (1.00000004) = 1.7371778928694496848392363956673867652098621469645354397627060605201847E-8
		x"0000000017371779241386000512000000000001145482042235960490901698081008", -- LUT(9) = log (1.000000004) = 1.7371779241386514646434499739319145482042235960490901698081007495768659E-9
		x"0000000001737177927265500000000000000000116070443631027431432640328547", -- LUT(10) = log (1.0000000004) = 1.7371779272655717251745637029904160704436310274314326403285426007813899E-10
		x"0000000000173717792757820005120000000000012915804974110630959916413016", -- LUT(11) = log (1.00000000004) = 1.7371779275782637520531820243490291580497411063095991641301789241946150E-11
		x"0000000000017371779276095000512000000000001585394037315649207411828745", -- LUT(12) = log (1.000000000004) = 1.7371779276095329547492989259941585394037315649207411828743800992112478E-12
		x"0000000000001737177927612600051200000000000188898708383124547867559775", -- LUT(13) = log (1.0000000000004) = 1.7371779276126598750189931668537888987083831245478675597769068803705788E-13
		x"0000000000000173717792761290005120000000000010313359098413228364926588", -- LUT(14) = log (1.00000000000004) = 1.7371779276129725670459634164467031335909841322836492658252404415865692E-14
		x"0000000000000017371779276130000256000000000001640690935060349023851518", -- LUT(15) = log (1.000000000000004) = 1.7371779276130038362486604496610640690935060349023851510772949189241865E-15
		x"0000000000000001737177927613000051200000000000150857763925583626037828", -- LUT(16) = log (1.0000000000000004) = 1.7371779276130069631689301530650508577639255836260378229344379240724406E-16
		x"0000000000000000173717792761300005120000000000017504358216923682346421", -- LUT(17) = log (1.00000000000000004) = 1.7371779276130072758609571234062750435821692368234642084675732156782286E-17
		x"0000000000000000017371779276130000000000000000001057172335056191511972", -- LUT(18) = log (1.000000000000000004) = 1.7371779276130073071301598204404057172335056191511979015318758479802509E-18
		x"0000000000000000001737177927613000000000000000000118867149334377554071", -- LUT(19) = log (1.0000000000000000004) = 1.7371779276130073102570800901438188671493343775540759218267435172142596E-19
		x"0000000000000000000173717792761300000000000000000016018296642420459603", -- LUT(20) = log (1.00000000000000000004) = 1.7371779276130073105697721171141601829664242045960647951065579857126789E-20
		x"0000000000000000000017371779276130000000000000000001943145563882568123", -- LUT(21) = log (1.000000000000000000004) = 1.7371779276130073106010413198111943145563882568122806931717831529057860E-21
		x"0000000000000000000001737177927613000000000000000000197727715467212724", -- LUT(22) = log (1.0000000000000000000004) = 1.7371779276130073106041682400808977277154672127290224530857028472718569E-22
		x"0000000000000000000000173717792761300000000000000000016806903137593385", -- LUT(23) = log (1.00000000000000000000004) = 1.7371779276130073106044809321078680690313759338276478307781688132253749E-23
		x"0000000000000000000000017371779276130000000000000000001651031629668148", -- LUT(24) = log (1.000000000000000000000004) = 1.7371779276130073106045122013105651031629668141925798805644261498106362E-24
		x"0000000000000000000000001737177927613000000000000000000134806576125909", -- LUT(25) = log (1.0000000000000000000000004) = 1.7371779276130073106045153282308348065761259023116237806632219908690862E-25
		x"0000000000000000000000000173717792761300000000000000000016177691744184", -- LUT(26) = log (1.00000000000000000000000004) = 1.7371779276130073106045156409228617769174418111243536776243032760489305E-26
		x"0000000000000000000000000017371779276130000000000000000001644739515734", -- LUT(27) = log (1.000000000000000000000000004) = 1.7371779276130073106045156721920644739515734020056349223899234215776549E-27
		x"0000000000000000000000000001737177927613000000000000000000184743654984", -- LUT(28) = log (1.0000000000000000000000000004) = 1.7371779276130073106045156753189847436549865610937631294171805563006347E-28
		x"0000000000000000000000000000173717792761300000000000000000017677062534", -- LUT(29) = log (1.00000000000000000000000000004) = 1.7371779276130073106045156756316767706253278770025759509454132209746338E-29
		x"0000000000000000000000000000017371779276130000000000000000001459733224", -- LUT(30) = log (1.000000000000000000000000000004) = 1.7371779276130073106045156756629459733223620085934572331064915569540507E-30
		x"0000000000000000000000000000001737177927613000000000000000000172893598", -- LUT(31) = log (1.0000000000000000000000000000004) = 1.7371779276130073106045156756660728935920654217525453613226819412471126E-31
		x"0000000000000000000000000000000173717792761300000000000000000018558567", -- LUT(32) = log (1.00000000000000000000000000000004) = 1.7371779276130073106045156756663855856190357630684541741443018051833699E-32
		x"0000000000000000000000000000000017371779276130000000000000000001168545", -- LUT(33) = log (1.000000000000000000000000000000004) = 1.7371779276130073106045156756664168548217327972000450554264637998320652E-33
		x"0000000000000000000000000000000001737177927613000000000000000000119986", -- LUT(34) = log (1.0000000000000000000000000000000004) = 1.7371779276130073106045156756664199817420025006132041435546799993794854E-34
		x"0000000000000000000000000000000000173717792761300000000000000000012024", -- LUT(35) = log (1.00000000000000000000000000000000004) = 1.7371779276130073106045156756664202944340294709545200523675016193350529E-35
		x"0000000000000000000000000000000000017371779276130000000000000000001202"); -- LUT(36) = log (1.000000000000000000000000000000000004) = 1.7371779276130073106045156756664202944340294709545200523675016193350529E-36

signal lut_LogShN5: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada0
		x"1760912590556800000000000000000122824319389827285873235194381791781200", -- LUT(1) = log (1.5) = 0.17609125905568124208128900853062228243193898272858732351943817917812096
		x"0211892990699380007680000000000014759155113790525527300230731328963749", -- LUT(2) = log (1.05) = 0.021189299069938072793505267123258475915511379052552730023073132896374403
		x"0021660617565076000256000000000001633815650632972011926373541806781619", -- LUT(3) = log (1.005) = 0.0021660617565076762304206377566908633815650632972011926373541806781611092
		x"0002170929722302000000000000000000133837444349518373528604405734453958", -- LUT(4) = log (1.0005) = 0.00021709297223020828191288375106682338374443495183735286044057344539553187
		x"0000217141812451550000000000000000011370670812814498785624291263197577", -- LUT(5) = log (1.00005) = 0.000021714181245155137172421675214706137067081281449878562429126319757005977
		x"0000021714669808533000768000000000001570878257409946699905137868615806", -- LUT(6) = log (1.000005) = 0.0000021714669808533308831621930838274570878257409946699905137868615805796951
		x"0000002171471866648300000000000000000175447233978551745997972670934195", -- LUT(7) = log (1.0000005) = 2.1714718666483377151571278999460754472339785517459979726709341906706011E-7
		x"0000000217147235522940000000000000000010938390090587995385342084310834", -- LUT(8) = log (1.00000005) = 2.1714723552294507099094395432311093839009058799538534208431083977367025E-8
		x"0000000021714724040875000256000000000001942178624117765985389455139813", -- LUT(9) = log (1.000000005) = 2.1714724040875781325606000937208942178624117765985389455139816328370259E-9
		x"0000000002171472408973300025600000000000110678243959366069409951126442", -- LUT(10) = log (1.0000000005) = 2.1714724089733910360575358440776106782439593660694099511264436608760878E-10
		x"0000000000217147240946190002560000000000012998737649442880279368602251", -- LUT(11) = log (1.00000000005) = 2.1714724094619723280195476764678299873764944288027936860225246918093730E-11
		x"0000000000021714724095108000512000000000001988676198334654162770405770", -- LUT(12) = log (1.000000000005) = 2.1714724095108304572318720423407988676198334654162770405776598533105943E-12
		x"0000000000002171472409515700051200000000000195626610408947838491761562", -- LUT(13) = log (1.0000000000005) = 2.1714724095157162701532657107544956266104089478384917615684286703025224E-13
		x"0000000000000217147240951620005120000000000012936162060187674995247933", -- LUT(14) = log (1.00000000000005) = 2.1714724095162048514454066899141293616206018767499524793820013234035099E-14
		x"0000000000000021714724095162000000000000000001753757731339964150883914", -- LUT(15) = log (1.000000000000005) = 2.1714724095162537095746208039532753757731339964150883915150616119884760E-15
		x"0000000000000002171472409516200076800000000000121803594962738122309425", -- LUT(16) = log (1.0000000000000005) = 2.1714724095162585953875422155184218035949627381223094201615105091033212E-16
		x"0000000000000000217147240951620007680000000000014876464121142799191156", -- LUT(17) = log (1.00000000000000005) = 2.1714724095162590839688343566765487646412114279919115649636746264634892E-17
		x"0000000000000000021714724095162000256000000000001775839284769551962627", -- LUT(18) = log (1.000000000000000005) = 2.1714724095162591328269635707923775839284769551962620528308318340922718E-18
		x"0000000000000000002171472409516200025600000000000160627089029914498938", -- LUT(19) = log (1.0000000000000000005) = 2.1714724095162591377127764922039606270890299144989314058243845286592757E-19
		x"0000000000000000000217147240951620002560000000000011893301740347449507", -- LUT(20) = log (1.00000000000000000005) = 2.1714724095162591382013577843451189330174034744950207445672811354198867E-20
		x"0000000000000000000021714724095162000256000000000001347636263640131357", -- LUT(21) = log (1.000000000000000000005) = 2.1714724095162591382502159135592347636263640131352879025364076824365528E-21
		x"0000000000000000000002171472409516200025600000000000146346687421298828", -- LUT(22) = log (1.0000000000000000000005) = 2.1714724095162591382551017264806463466874212988257212005743291074745930E-22
		x"0000000000000000000000217147240951620002560000000000018750499352863979", -- LUT(23) = log (1.00000000000000000000005) = 2.1714724095162591382555903077727875049935286397130285962005313980832338E-23
		x"0000000000000000000000021714724095162000256000000000001016208241393895", -- LUT(24) = log (1.000000000000000000000005) = 2.1714724095162591382556391659020016208241393899249419764213757286855477E-24
		x"0000000000000000000000002171472409516200025600000000000123032407200464", -- LUT(25) = log (1.0000000000000000000000005) = 2.1714724095162591382556440517149230324072004651073651408500424027612540E-25
		x"0000000000000000000000000217147240951620002560000000000011517356550653", -- LUT(26) = log (1.00000000000000000000000005) = 2.1714724095162591382556445402962151735655065726272197755569748925789794E-26
		x"0000000000000000000000000021714724095162000256000000000001443876813372", -- LUT(27) = log (1.000000000000000000000000005) = 2.1714724095162591382556445891543443876813371833792213622103087997848535E-27
		x"0000000000000000000000000002171472409516200025600000000000157309092921", -- LUT(28) = log (1.0000000000000000000000000005) = 2.1714724095162591382556445940401573090929202444544216821074685970876819E-28
		x"0000000000000000000000000000217147240951620002560000000000013860123400", -- LUT(29) = log (1.00000000000000000000000000005) = 2.1714724095162591382556445945287386012340785505619417157095028408837872E-29
		x"0000000000000000000000000000021714724095162000256000000000001967304480", -- LUT(30) = log (1.000000000000000000000000000005) = 2.1714724095162591382556445945775967304481943811726937190858294479040559E-30
		x"0000000000000000000000000000002171472409516200025600000000000182543367", -- LUT(31) = log (1.0000000000000000000000000000005) = 2.1714724095162591382556445945824825433696059642337689194236233404324894E-31
		x"0000000000000000000000000000000217147240951620002560000000000017112465", -- LUT(32) = log (1.00000000000000000000000000000005) = 2.1714724095162591382556445945829711246617471225398764394574043420035968E-32
		x"0000000000000000000000000000000021714724095162000256000000000001199825", -- LUT(33) = log (1.000000000000000000000000000000005) = 2.1714724095162591382556445945830199827909612383704871914607824582838902E-33
		x"0000000000000000000000000000000002171472409516200025600000000000124864", -- LUT(34) = log (1.0000000000000000000000000000000005) = 2.1714724095162591382556445945830248686038826499535482666611202700731513E-34
		x"0000000000000000000000000000000000217147240951620002560000000000012533", -- LUT(35) = log (1.00000000000000000000000000000000005) = 2.1714724095162591382556445945830253571851747911118543741811540512536898E-35
		x"0000000000000000000000000000000000021714724095162000256000000000001253"); -- LUT(36) = log (1.000000000000000000000000000000000005) = 2.1714724095162591382556445945830253571851747911118543741811540512536898E-36

signal lut_LogShN4: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2041199826559200000000000000000121070727595258484341652417098445084320", -- LUT(1) = log (1.6) = 0.20411998265592478085495557889797210707275952584843416524170984450843276
		x"0253058652647700007680000000000016194636922827570463219045304169023330", -- LUT(2) = log (1.06) = 0.025305865264770240846731186351749619463692282757046321904530416902333994
		x"0025979807199085000000000000000001817743691929947498513731263267939608", -- LUT(3) = log (1.006) = 0.0025979807199085923119629850040210817743691929947498513731263267939609060
		x"0002604985473903400076800000000000190107995813225361469363224218313447", -- LUT(4) = log (1.0006) = 0.00026049854739034681785461091743713901079958132253614693632242183134479412
		x"0000260568872153950002560000000000013603269126525260588336231493027868", -- LUT(5) = log (1.00006) = 0.000026056887215395479456228829083273360326912652526058833623149302786684559
		x"0000026057590741501000512000000000001785317512066118325462073039515087", -- LUT(6) = log (1.000006) = 0.0000026057590741501057693601731995175785317512066118325462073039515082024391
		x"0000002605766109689700025600000000000175719412067329744741644439916436", -- LUT(7) = log (1.0000006) = 2.6057661096897562319397427381882757194120673297447416444399164380100951E-7
		x"0000000260576681324650002560000000000010167075837645628087129931819085", -- LUT(8) = log (1.00000006) = 2.6057668132465073502415735283042016707583764562808712993181908973059563E-8
		x"0000000026057668836022000000000000000001300829099554354160179395952374", -- LUT(9) = log (1.000000006) = 2.6057668836022103229174431721020300829099554354160179395952376904460728E-9
		x"0000000002605766890637700076800000000000128343556193593944897661103985", -- LUT(10) = log (1.0000000006) = 2.6057668906377808987936122505572283435561935939448976611039831934307910E-10
		x"0000000000260576689134130005120000000000018999010835134878083074812985", -- LUT(11) = log (1.00000000006) = 2.6057668913413379591673151047919899901083513487808307481298879152458436E-11
		x"0000000000026057668914116000512000000000001070666460618886446848654345", -- LUT(12) = log (1.000000000006) = 2.6057668914116936652325462498046070666460618886446848654349723368812723E-12
		x"0000000000002605766891418700025600000000000185431912936642350105051355", -- LUT(13) = log (1.0000000000006) = 2.6057668914187292358393479729018854319129366423501050513507951413665434E-13
		x"0000000000000260576689141940007680000000000017356026424949358317797455", -- LUT(14) = log (1.00000000000006) = 2.6057668914194327929000309312975735602642494935831779745872234483222515E-14
		x"0000000000000026057668914195000256000000000001019761428755268099872434", -- LUT(15) = log (1.000000000000006) = 2.6057668914195031486060992549980019761428755268099872430496970547346806E-15
		x"0000000000000002605766891419500076800000000000153413761298326108048663", -- LUT(16) = log (1.0000000000000006) = 2.6057668914195101841767060876466534137612983261080486674570786834371329E-16
		x"0000000000000000260576689141950007680000000000010464348344633324610292", -- LUT(17) = log (1.00000000000000006) = 2.6057668914195108877337667709143046434834463332461029604113412003063937E-17
		x"0000000000000000026057668914195000512000000000001976273152641913572392", -- LUT(18) = log (1.000000000000000006) = 2.6057668914195109580894728392410976273152641913572393655574466198711641E-18
		x"0000000000000000002605766891419500051200000000000177204307042007742451", -- LUT(19) = log (1.0000000000000000006) = 2.6057668914195109651250434460737772043070420077424515643249094980318901E-19
		x"0000000000000000000260576689141950005120000000000014516479230574968671", -- LUT(20) = log (1.00000000000000000006) = 2.6057668914195109658286005067570451647923057496867138950326786547545908E-20
		x"0000000000000000000026057668914195000512000000000001719608686929834842", -- LUT(21) = log (1.000000000000000000006) = 2.6057668914195109658989562128253719608686929834841975393370142934614718E-21
		x"0000000000000000000002605766891419500051200000000000104640476610315454", -- LUT(22) = log (1.0000000000000000000006) = 2.6057668914195109659059917834322046404766103154599764778799086930568515E-22
		x"0000000000000000000000260576689141950005120000000000018790843740483478", -- LUT(23) = log (1.00000000000000000000006) = 2.6057668914195109659066953404928879084374048347435146774753228666221307E-23
		x"0000000000000000000000026057668914195000512000000000001562352334843147", -- LUT(24) = log (1.000000000000000000000006) = 2.6057668914195109659067656961989562352334843145327281004922755314399646E-24
		x"0000000000000000000000002605766891419500051200000000000163067913092267", -- LUT(25) = log (1.0000000000000000000000006) = 2.6057668914195109659067727317695630679130922627902580388245449103964863E-25
		x"0000000000000000000000000260576689141950005120000000000012375118105307", -- LUT(26) = log (1.00000000000000000000000006) = 2.6057668914195109659067734353266237511810530576187971186180775894168859E-26
		x"0000000000000000000000000026057668914195000512000000000001298195078497", -- LUT(27) = log (1.000000000000000000000000006) = 2.6057668914195109659067735056823298195078491371016788874570339147301734E-27
		x"0000000000000000000000000002605766891419500051200000000000100426340526", -- LUT(28) = log (1.0000000000000000000000000006) = 2.6057668914195109659067735127179004263405287450499673429495255778356146E-28
		x"0000000000000000000000000000260576689141950005120000000000015748702375", -- LUT(29) = log (1.00000000000000000000000000006) = 2.6057668914195109659067735134214574870237967058447961912848607044518998E-29
		x"0000000000000000000000000000026057668914195000512000000000001131930923", -- LUT(30) = log (1.000000000000000000000000000006) = 2.6057668914195109659067735134918131930921235019242790761462550767165858E-30
		x"0000000000000000000000000000002605766891419500051200000000000148763690", -- LUT(31) = log (1.0000000000000000000000000000006) = 2.6057668914195109659067735134988487636989561815322273646326731225390850E-31
		x"0000000000000000000000000000000260576689141950005120000000000015232072", -- LUT(32) = log (1.00000000000000000000000000000006) = 2.6057668914195109659067735134995523207596394494930221934813177132072952E-32
		x"0000000000000000000000000000000026057668914195000512000000000001226761", -- LUT(33) = log (1.000000000000000000000000000000006) = 2.6057668914195109659067735134996226764657077762891016763661822001349758E-33
		x"0000000000000000000000000000000002605766891419500051200000000000129718", -- LUT(34) = log (1.0000000000000000000000000000000006) = 2.6057668914195109659067735134996297120363146089687096246546686491063525E-34
		x"0000000000000000000000000000000000260576689141950005120000000000013040", -- LUT(35) = log (1.00000000000000000000000000000000006) = 2.6057668914195109659067735134996304155933752922366704194835172940062762E-35
		x"0000000000000000000000000000000000026057668914195000512000000000001304"); -- LUT(36) = log (1.000000000000000000000000000000000006) = 2.6057668914195109659067735134996304155933752922366704194835172940062762E-36

signal lut_LogShN3: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2304489213782700076800000000000170300075673784250463973803684823446940", -- LUT(1) = log (1.7) = 0.23044892137827392854016989432833703000756737842504639738036848234469406
		x"0293837776852090007680000000000016461268168916340193519816620084607712", -- LUT(2) = log (1.07) = 0.029383777685209640834541239461435646126816891634019351981662008460771940
		x"0030294705536180000512000000000001106466317386894353795009218244829763", -- LUT(3) = log (1.007) = 0.0030294705536180071693257673841859106466317386894353795009218244829766464
		x"0003038997848124900000000000000000144183182228888561508963181665084194", -- LUT(4) = log (1.0007) = 0.00030389978481249181051766773638472441831822288885615089631816650841904241
		x"0000303995497613980000000000000000019256695912333182293488937204796115", -- LUT(5) = log (1.00007) = 0.000030399549761398694026220679023281925669591233318229348893720479611201115
		x"0000030400507331576000256000000000001937458283326137859440297095332826", -- LUT(6) = log (1.000007) = 0.0000030400507331576102389685938385813937458283326137859440297095332822755125
		x"0000003040060309301700051200000000000167101385693171650278081171046767", -- LUT(7) = log (1.0000007) = 3.0400603093017786736878822882945671013856931716502780811710467620915983E-7
		x"0000000304006126692060007680000000000011586635341666788797292950894478", -- LUT(8) = log (1.00000007) = 3.0400612669206196926945203998207158663534166678879729295089447889260909E-8
		x"0000000030400613626825000256000000000001080547935809934934811381154279", -- LUT(9) = log (1.000000007) = 3.0400613626825480365825681585501080547935809934934811381154272700479085E-9
		x"0000000003040061372258700000000000000000102385046444157146590192654448", -- LUT(10) = log (1.0000000007) = 3.0400613722587413133914788120530023850464441571465901926544471003248430E-10
		x"0000000000304006137321630002560000000000017548489294087423498480202161", -- LUT(11) = log (1.00000000007) = 3.0400613732163606454965711682178754848929408742349848020216741125759402E-11
		x"0000000000030400613733121000768000000000001469286543542342154439585444", -- LUT(12) = log (1.000000000007) = 3.0400613733121225787513224169745469286543542342154439585443370392063612E-12
		x"0000000000003040061373321600051200000000000147952666671043202494392325", -- LUT(13) = log (1.0000000000007) = 3.0400613733216987720772399619818479526666710432024943923216583293337840E-13
		x"0000000000000304006137332260007680000000000019462590256301659564872956", -- LUT(14) = log (1.00000000000007) = 3.0400613733226563914098361406838946259025630165956487295034331493131026E-14
		x"0000000000000030400613733227000512000000000001124591665371154106660607", -- LUT(15) = log (1.000000000000007) = 3.0400613733227521533430958027961124591665371154106660607118830966205115E-15
		x"0000000000000003040061373322700025600000000000154374152570412605476868", -- LUT(16) = log (1.0000000000000007) = 3.0400613733227617295364217694497543741525704126054768694967134847582125E-16
		x"0000000000000000304006137332270007680000000000014276696777033323638953", -- LUT(17) = log (1.00000000000000007) = 3.0400613733227626871557543661195427669677703332363895933184539132192355E-17
		x"0000000000000000030400613733227000768000000000001658482624562914406332", -- LUT(18) = log (1.000000000000000007) = 3.0400613733227627829176876257865658482624562914406334806822601403428280E-18
		x"0000000000000000003040061373322700076800000000000168598812056546922701", -- LUT(19) = log (1.0000000000000000007) = 3.0400613733227627924938809517532685988120565469227014338670092858076277E-19
		x"0000000000000000000304006137332270007680000000000013887829121788906751", -- LUT(20) = log (1.00000000000000000007) = 3.0400613733227627934515002843499388782912178890675248968682664377826717E-20
		x"0000000000000000000030400613733227000768000000000001059062833760364472", -- LUT(21) = log (1.000000000000000000007) = 3.0400613733227627935472622176096059062833760364479734100772582739066627E-21
		x"0000000000000000000003040061373322700076800000000000172609083034271313", -- LUT(22) = log (1.0000000000000000000007) = 3.0400613733227627935568384109355726090830342713176779230674781570268789E-22
		x"0000000000000000000000304006137332270007680000000000016927936300451904", -- LUT(23) = log (1.00000000000000000000007) = 3.0400613733227627935577960302681692793630045190059649709831935843722773E-23
		x"0000000000000000000000030400613733227000768000000000001289463910015885", -- LUT(24) = log (1.000000000000000000000007) = 3.0400613733227627935578917922014289463910015880168068417409320617291892E-24
		x"0000000000000000000000003040061373322700076800000000000154913093801296", -- LUT(25) = log (1.0000000000000000000000007) = 3.0400613733227627935579013683947549130938012953603111604763675788113361E-25
		x"0000000000000000000000000304006137332270007680000000000018750976408127", -- LUT(26) = log (1.00000000000000000000000007) = 3.0400613733227627935579023260140875097640812660990857936665077472130156E-26
		x"0000000000000000000000000030400613733227000768000000000001207694311095", -- LUT(27) = log (1.000000000000000000000000007) = 3.0400613733227627935579024217760207694311092631730074989986877302201182E-27
		x"0000000000000000000000000003040061373322700076800000000000114095397814", -- LUT(28) = log (1.0000000000000000000000000007) = 3.0400613733227627935579024313522140953978120628804001119520373881824978E-28
		x"0000000000000000000000000000304006137332270007680000000000013342799443", -- LUT(29) = log (1.00000000000000000000000000007) = 3.0400613733227627935579024323098334279944823428511393776715736705753525E-29
		x"0000000000000000000000000000030400613733227000768000000000001953612543", -- LUT(30) = log (1.000000000000000000000000000007) = 3.0400613733227627935579024324055953612541493708482133042877693119806041E-30
		x"0000000000000000000000000000003040061373322700076800000000000171554588", -- LUT(31) = log (1.0000000000000000000000000000007) = 3.0400613733227627935579024324151715545801160736479206969498312962527889E-31
		x"0000000000000000000000000000000304006137332270007680000000000012917399", -- LUT(32) = log (1.00000000000000000000000000000007) = 3.0400613733227627935579024324161291739127127439278914362160419188813240E-32
		x"0000000000000000000000000000000030400613733227000768000000000001249355", -- LUT(33) = log (1.000000000000000000000000000000007) = 3.0400613733227627935579024324162249358459724109558885101426630253861907E-33
		x"0000000000000000000000000000000003040061373322700076800000000000134514", -- LUT(34) = log (1.0000000000000000000000000000000007) = 3.0400613733227627935579024324162345120392983776586882175353251364790975E-34
		x"0000000000000000000000000000000000304006137332270007680000000000013543", -- LUT(35) = log (1.00000000000000000000000000000000007) = 3.0400613733227627935579024324162354696586309743289681882745913475928123E-35
		x"0000000000000000000000000000000000030400613733227000768000000000001354"); -- LUT(36) = log (1.000000000000000000000000000000000007) = 3.0400613733227627935579024324162354696586309743289681882745913475928123E-36

signal lut_LogShN2: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2552725051033000076800000000000136451684476098435002709701587417375660", -- LUT(1) = log (1.8) = 0.25527250510330606980379470123472364516844760984350027097015874173756649
		x"0334237554869490002560000000000019811367663554963046771104518431699035", -- LUT(2) = log (1.08) = 0.033423755486949702312561499214331981136766355496304677110451843169903837
		x"0034605321095064000512000000000001189565896505537913014050760788371445", -- LUT(3) = log (1.008) = 0.0034605321095064861572276440008389189565896505537913014050760788371445026
		x"0003472966853635400076800000000000131845603406855766932484444966633035", -- LUT(4) = log (1.0008) = 0.00034729668536354068770569300355701318456034068557669324844449666330305433
		x"0000347421688840330002560000000000019207216874281586059046883252658513", -- LUT(5) = log (1.00008) = 0.000034742168884033200493502377533561920721687428158605904688325265851489058
		x"0000034743419578767000512000000000001722989729673547644029504139573582", -- LUT(6) = log (1.000008) = 0.0000034743419578767128640139981982054722989729673547644029504139573588112687
		x"0000003474354465484400025600000000000170094483230281108248532617587241", -- LUT(7) = log (1.0000008) = 3.4743544654844137262742471526562700944832302811082485326175872406141605E-7
		x"0000000347435571625170000000000000000013817570546789709054114330912102", -- LUT(8) = log (1.00000008) = 3.4743557162517878241271596009484381757054678970905411433091210037269144E-8
		x"0000000034743558413285000512000000000001472160789083532224132159169319", -- LUT(9) = log (1.000000008) = 3.4743558413285912744245639999341472160789083532224132159169313812007575E-9
		x"0000000003474355853836200076800000000000160354495655831327214401281878", -- LUT(10) = log (1.0000000008) = 3.4743558538362722798598214181860603544956558313272144012818766245188488E-10
		x"0000000000347435585508700007680000000000015018461100121902961823850020", -- LUT(11) = log (1.00000000008) = 3.4743558550870403870074027256418501846110012190296182385002100765274322E-11
		x"0000000000034743558552121000768000000000001822432108810103810610604905", -- LUT(12) = log (1.000000000008) = 3.4743558552121171977882014124395822432108810103810610604901214372805351E-12
		x"0000000000003474355855224600076800000000000172826919711218624033490554", -- LUT(13) = log (1.0000000000008) = 3.4743558552246248788669416866802728269197112186240334905533028938205856E-13
		x"0000000000000347435585522580002560000000000015145491617587383279630333", -- LUT(14) = log (1.00000000000008) = 3.4743558552258756469748223181599514549161758738327963033075749065134465E-14
		x"0000000000000034743558552260000000000000000001754138079252489349423082", -- LUT(15) = log (1.000000000000008) = 3.4743558552260007237856104473484754138079252489349423081128531596023001E-15
		x"0000000000000003474355855226000025600000000000133370658417062634209561", -- LUT(16) = log (1.0000000000000008) = 3.4743558552260132314666892609277333706584170626342095640645664460388304E-16
		x"0000000000000000347435585522600007680000000000016322195307980861312008", -- LUT(17) = log (1.00000000000000008) = 3.4743558552260144822347971422922632219530798086131200564260023217039677E-17
		x"0000000000000000034743558552260000000000000000001822476386422192529487", -- LUT(18) = log (1.000000000000000008) = 3.4743558552260146073116079304287822476386422192529480365700454391136525E-18
		x"0000000000000000003474355855226000000000000000000134810612759421677747", -- LUT(19) = log (1.0000000000000000008) = 3.4743558552260146198192890092424348106127594216777460509867689855705937E-19
		x"0000000000000000000347435585522600000000000000000010007351422675153386", -- LUT(20) = log (1.00000000000000000008) = 3.4743558552260146210700571171238000735142267515338344004395577728031184E-20
		x"0000000000000000000034743558552260000000000000000001365998704140406155", -- LUT(21) = log (1.000000000000000000008) = 3.4743558552260146211951339279119365998704140406155793212607949090924788E-21
		x"0000000000000000000003474355855226000000000000000000150252506693175084", -- LUT(22) = log (1.0000000000000000000008) = 3.4743558552260146212076416089907502525066931750847151742020740523903162E-22
		x"0000000000000000000000347435585522600000000000000000013161777032769253", -- LUT(23) = log (1.00000000000000000000008) = 3.4743558552260146212088923770986316177703276925872383731047939168638822E-23
		x"0000000000000000000000034743558552260000000000000000001197542966912102", -- LUT(24) = log (1.000000000000000000000008) = 3.4743558552260146212090174539094197542966912103780467891311518232085237E-24
		x"0000000000000000000000003474355855226000000000000000000198567949327561", -- LUT(25) = log (1.0000000000000000000000008) = 3.4743558552260146212090299615904985679493275628175331916951484730423565E-25
		x"0000000000000000000000000347435585522600000000000000000010644931459110", -- LUT(26) = log (1.00000000000000000000000008) = 3.4743558552260146212090312123586064493145911980680858875611617466177339E-26
		x"0000000000000000000000000034743558552260000000000000000001172374511177", -- LUT(27) = log (1.000000000000000000000000008) = 3.4743558552260146212090313374354172374511175615932071977038592100611916E-27
		x"0000000000000000000000000003474355855226000000000000000000198316264776", -- LUT(28) = log (1.0000000000000000000000000008) = 3.4743558552260146212090313499430983162647701979457199891236899177663966E-28
		x"0000000000000000000000000000347435585522600000000000000000016642414615", -- LUT(29) = log (1.00000000000000000000000000008) = 3.4743558552260146212090313511938664241461354615809712748697285981505256E-29
		x"0000000000000000000000000000034743558552260000000000000000001432349344", -- LUT(30) = log (1.000000000000000000000000000008) = 3.4743558552260146212090313513189432349342719879444964035103730222850746E-30
		x"0000000000000000000000000000003474355855226000000000000000000150916013", -- LUT(31) = log (1.0000000000000000000000000000008) = 3.4743558552260146212090313513314509160130856405808489163750978702594909E-31
		x"0000000000000000000000000000000347435585522600000000000000000010168412", -- LUT(32) = log (1.00000000000000000000000000000008) = 3.4743558552260146212090313513327016841209670058444841676615769591125421E-32
		x"0000000000000000000000000000000034743558552260000000000000000001267601", -- LUT(33) = log (1.000000000000000000000000000000008) = 3.4743558552260146212090313513328267609317551423708476927902249340384034E-33
		x"0000000000000000000000000000000003474355855226000000000000000000139269", -- LUT(34) = log (1.0000000000000000000000000000000008) = 3.4743558552260146212090313513328392686128339560234840453030897321913950E-34
		x"0000000000000000000000000000000000347435585522600000000000000000014058", -- LUT(35) = log (1.00000000000000000000000000000000008) = 3.4743558552260146212090313513328405193809418373887476805543762120132983E-35
		x"0000000000000000000000000000000000034743558552260000000000000000001405"); -- LUT(36) = log (1.000000000000000000000000000000000008) = 3.4743558552260146212090313513328405193809418373887476805543762120132983E-36

signal lut_LogShN1: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"2787536009528200000000000000000193179511293373944975989068188687077500", -- LUT(1) = log (1.9) = 0.27875360095282896153633347575692931795112933739449759890681886870775084
		x"0374264979406230000000000000000012866422045228279836821104005352703150", -- LUT(2) = log (1.09) = 0.037426497940623635200513307613875286642204522827983682110400535270315801
		x"0038911662369105000000000000000001655201956525526009846382285243403377", -- LUT(3) = log (1.009) = 0.0038911662369105217152813165095588655201956525526009846382285243403377898
		x"0003906892499101300076800000000000177117353304961609395099081154215706", -- LUT(4) = log (1.0009) = 0.00039068924991013102886422325456872771173533049616093950990811542157087625
		x"0000390847445841670002560000000000018620649738205286721679085600295386", -- LUT(5) = log (1.00009) = 0.000039084744584167392418805024884522862064973820528672167908560029538579932
		x"0000039086327483082000000000000000001391142079074510492256220353603875", -- LUT(6) = log (1.000009) = 0.0000039086327483082822139172355443443391142079074510492256220353603872872196
		x"0000003908648578237600051200000000000120129943352801981548597095287414", -- LUT(7) = log (1.0000009) = 3.9086485782376700755689321740694201299433528019815485970952874117444642E-7
		x"0000000390865016124000002560000000000019299892405193409790258911024413", -- LUT(8) = log (1.00000009) = 3.9086501612400118313983679690889929989240519340979025891102441904109279E-8
		x"0000000039086503195403000256000000000001998308735181253221841864747612", -- LUT(9) = log (1.000000009) = 3.9086503195403400373120196405173998308735181253221841864747610661621882E-9
		x"0000000003908650335370300076800000000000124036800650028456709883035251", -- LUT(10) = log (1.0000000009) = 3.9086503353703737982073259585749240368006500284567098830352564584361153E-10
		x"0000000000390865033695330007680000000000017519637637990713285701050625", -- LUT(11) = log (1.00000000009) = 3.9086503369533771836998966359602751963763799071328570105062129289720063E-11
		x"0000000000039086503371116000000000000000001767972760458340474934189089", -- LUT(12) = log (1.000000000009) = 3.9086503371116775223431841047886767972760458340474934189083802899778119E-12
		x"0000000000003908650337127500051200000000000149692717550469951683837298", -- LUT(13) = log (1.0000000000009) = 3.9086503371275075562084531556830496927175504699516838372994026827053774E-13
		x"0000000000000390865033712900005120000000000010294368571888757316083637", -- LUT(14) = log (1.00000000000009) = 3.9086503371290905595949894638126029436857188875731608363952420228844874E-14
		x"0000000000000039086503371292000512000000000001594290308464114948665576", -- LUT(15) = log (1.000000000000009) = 3.9086503371292488599336431886559594290308464114948665574444026612025644E-15
		x"0000000000000003908650337129200076800000000000199089168476341211256525", -- LUT(16) = log (1.0000000000000009) = 3.9086503371292646899675085620805990891684763412112565220533695965814975E-16
		x"0000000000000000390865033712920005120000000000016609529827114002664034", -- LUT(17) = log (1.00000000000000009) = 3.9086503371292662729708950994324660952982711400266403367080845627523069E-17
		x"0000000000000000039086503371292000256000000000001468263124109386006863", -- LUT(18) = log (1.000000000000000009) = 3.9086503371292664312712337531677468263124109386006866689798086683705157E-18
		x"0000000000000000003908650337129200025600000000000175839717836521645652", -- LUT(19) = log (1.0000000000000000009) = 3.9086503371292664471012676185412758397178365216456504522176679240134738E-19
		x"0000000000000000000390865033712920002560000000000012875046141919598201", -- LUT(20) = log (1.00000000000000000009) = 3.9086503371292664486842710050786287504614191959820230561120633423480286E-20
		x"0000000000000000000039086503371292000256000000000001640416298078645759", -- LUT(21) = log (1.000000000000000000009) = 3.9086503371292664488425713437323640416298078645759790793912794817335061E-21
		x"0000000000000000000003908650337129200025600000000000137570747587035448", -- LUT(22) = log (1.0000000000000000000009) = 3.9086503371292664488584013775977375707475870354469778693487329321501984E-22
		x"0000000000000000000000390865033712920002560000000000017492365937435557", -- LUT(23) = log (1.00000000000000000000009) = 3.9086503371292664488599843809842749236593743555741937802207742296271517E-23
		x"0000000000000000000000039086503371292000256000000000001286589505531816", -- LUT(24) = log (1.000000000000000000000009) = 3.9086503371292664488601426813229286589505531816173165316267413195332704E-24
		x"0000000000000000000000003908650337129200025600000000000194032479671065", -- LUT(25) = log (1.0000000000000000000000009) = 3.9086503371292664488601585113567940324796710651619328183705256581261006E-25
		x"0000000000000000000000000390865033712920002560000000000018056983258284", -- LUT(26) = log (1.00000000000000000000000009) = 3.9086503371292664488601600943601805698325828535257974871609359682814064E-26
		x"0000000000000000000000000039086503371292000256000000000001192235678743", -- LUT(27) = log (1.000000000000000000000000009) = 3.9086503371292664488601602526605192235678740323622779844411373180598972E-27
		x"0000000000000000000000000003908650337129200025600000000000153088941402", -- LUT(28) = log (1.0000000000000000000000000009) = 3.9086503371292664488601602684905530889414031502459269744731690562253759E-28
		x"0000000000000000000000000000390865033712920002560000000000015647547871", -- LUT(29) = log (1.00000000000000000000000000009) = 3.9086503371292664488601602700735564754787560620342918828794123460738001E-29
		x"0000000000000000000000000000039086503371292000256000000000001568141328", -- LUT(30) = log (1.000000000000000000000000000009) = 3.9086503371292664488601602702318568141324913532131283738140670762189613E-30
		x"0000000000000000000000000000003908650337129200025600000000000186847997", -- LUT(31) = log (1.0000000000000000000000000000009) = 3.9086503371292664488601602702476868479978648823310120229084728532450806E-31
		x"0000000000000000000000000000000390865033712920002560000000000016985136", -- LUT(32) = log (1.00000000000000000000000000000009) = 3.9086503371292664488601602702492698513844022352428003878179228339878085E-32
		x"0000000000000000000000000000000039086503371292000256000000000001281515", -- LUT(33) = log (1.000000000000000000000000000000009) = 3.9086503371292664488601602702494281517230559705339792243088679260924825E-33
		x"0000000000000000000000000000000003908650337129200025600000000000143984", -- LUT(34) = log (1.0000000000000000000000000000000009) = 3.9086503371292664488601602702494439817569213440630971079579624362432539E-34
		x"0000000000000000000000000000000000390865033712920002560000000000014553", -- LUT(35) = log (1.00000000000000000000000000000000009) = 3.9086503371292664488601602702494455647603078814160088963228718872677341E-35
		x"0000000000000000000000000000000000039086503371292000256000000000001455"); -- LUT(36) = log (1.000000000000000000000000000000000009) = 3.9086503371292664488601602702494455647603078814160088963228718872677341E-36

signal lut_LogShN0: mlut_LogShN := (
		x"0000000000000000000000000000000000000000000000000000000000000000000000", -- LUT(0), No usada
		x"3010299956639800051200000000000130267681898814621085413104274611271080", -- LUT(1) = log (2.0) = 0.30102999566398119521373889472449302676818988146210854131042746112710819
		x"0413926851582250005120000000000012417067021904664530945965390186797530", -- LUT(2) = log (1.10) = 0.041392685158225040750199971243024241706702190466453094596539018679753032
		x"0043213737826425000512000000000001132192893552064525914058186369484480", -- LUT(3) = log (1.010) = 0.0043213737826425742751881782229379132192893552064525914058186369484480104
		x"0004340774793186400076800000000000160200037751774867729013649473955590", -- LUT(4) = log (1.0010) = 0.00043407747931864066892138777798886602000377517748677290136494739555956377
		x"0000434272768626690002560000000000011310979627758925307732464042115847", -- LUT(5) = log (1.00010) = 0.000043427276862669637313527585098268131097962775892530773246404211584759011
		x"0000043429231044531000512000000000001839724439448249094541443880968626", -- LUT(6) = log (1.000010) = 0.0000043429231044531868554934716343971839724439448249094541443880968627435425
		x"0000004342942647561500000000000000000170416841361667145121612010092065", -- LUT(7) = log (1.0000010) = 4.3429426475615564074394264367770704168413616671451216120100920600646163E-7
		x"0000000434294460188520000000000000000014716184534126294027719584836884", -- LUT(8) = log (1.00000010) = 4.3429446018852918013670197358779471618453412629402771958483688371187471E-8
		x"0000000043429447973177000256000000000001513552500188036530684122042803", -- LUT(9) = log (1.000000010) = 4.3429447973177943261135240219573513552500188036530684122042800710352334E-9
		x"0000000004342944816861000051200000000000109449975167103574888128566602", -- LUT(10) = log (1.0000000010) = 4.3429448168610458684426783228355094499751671035748881285666077943342844E-10
		x"0000000000434294481881530002560000000000010902153603387684726625081271", -- LUT(11) = log (1.00000000010) = 4.3429448188153710355741397580695090215360338768472662508127253947631500E-11
		x"0000000000043429448190108000512000000000001943752044854307845718560522", -- LUT(12) = log (1.000000000010) = 4.3429448190108035524162713626107943752044854307845718560521428168814761E-12
		x"0000000000004342944819030300000000000000000168188103076331630995751303", -- LUT(13) = log (1.0000000000010) = 4.3429448190303468041017743776760681881030763316309957513017772960244133E-13
		x"0000000000000434294481903230002560000000000010798859182027432839105044", -- LUT(14) = log (1.00000000000010) = 4.3429448190323011292703375777287079885918202743283910504849072998679919E-14
		x"0000000000000043429448190324000512000000000001330937991070845967224895", -- LUT(15) = log (1.000000000000010) = 4.3429448190324965617871940267194330937991070845967224894788994375775741E-15
		x"0000000000000004342944819032500000000000000000160215572386313351021740", -- LUT(16) = log (1.0000000000000010) = 4.3429448190325161050388796729083602155723863133510217474644354630612721E-16
		x"0000000000000000434294481903250005120000000000015147386224070812729380", -- LUT(17) = log (1.00000000000000010) = 4.3429448190325180593640482375401514738622407081272938153719073538458377E-17
		x"0000000000000000043429448190325000512000000000001595851523514132903530", -- LUT(18) = log (1.000000000000000010) = 4.3429448190325182547965650940034595851523514132903530110647890888807852E-18
		x"0000000000000000004342944819032500051200000000000191686135973736464476", -- LUT(19) = log (1.0000000000000000010) = 4.3429448190325182743398167796497916861359737364644796740905796609375344E-19
		x"0000000000000000000434294481903250005120000000000012490913288208130847", -- LUT(20) = log (1.00000000000000000010) = 4.3429448190325182762941419482144249091328820813084715142512912231826086E-20
		x"0000000000000000000043429448190325000512000000000001882315615583769188", -- LUT(21) = log (1.000000000000000000010) = 4.3429448190325182764895744650708882315615583769181364909723672719385639E-21
		x"0000000000000000000004342944819032500051200000000000134563805715861099", -- LUT(22) = log (1.0000000000000000000010) = 4.3429448190325182765091177167565345638057158610903556465724913493069550E-22
		x"0000000000000000000000434294481903250005120000000000019919703014450809", -- LUT(23) = log (1.00000000000000000000010) = 4.3429448190325182765110720419250991970301445080536900887117848881922896E-23
		x"0000000000000000000000043429448190325000512000000000001556603525875019", -- LUT(24) = log (1.000000000000000000000010) = 4.3429448190325182765112674744419556603525875017354846581915070543587315E-24
		x"0000000000000000000000004342944819032500051200000000000141306684831809", -- LUT(25) = log (1.0000000000000000000000010) = 4.3429448190325182765112870176936413066848318023935187263921371990991212E-25
		x"0000000000000000000000000434294481903250005120000000000010987131805628", -- LUT(26) = log (1.00000000000000000000000010) = 4.3429448190325182765112889720188098713180562324722206793247267928543986E-26
		x"0000000000000000000000000043429448190325000512000000000001267277813787", -- LUT(27) = log (1.000000000000000000000000010) = 4.3429448190325182765112891674513267277813786754802198600791110180227388E-27
		x"0000000000000000000000000004342944819032500051200000000000178413427716", -- LUT(28) = log (1.0000000000000000000000000010) = 4.3429448190325182765112891869945784134277109197810210680091606931975009E-28
		x"0000000000000000000000000000434294481903250005120000000000010358199235", -- LUT(29) = log (1.00000000000000000000000000010) = 4.3429448190325182765112891889489035819923441442111012017007117732415564E-29
		x"0000000000000000000000000000043429448190325000512000000000001360988484", -- LUT(30) = log (1.000000000000000000000000000010) = 4.3429448190325182765112891891443360988488074666541092151988523423712277E-30
		x"0000000000000000000000000000004342944819032500051200000000000179350533", -- LUT(31) = log (1.0000000000000000000000000000010) = 4.3429448190325182765112891891638793505344537988984100165499562538954475E-31
		x"0000000000000000000000000000000434294481903250005120000000000013367572", -- LUT(32) = log (1.00000000000000000000000000000010) = 4.3429448190325182765112891891658336757030184321228400966850795435939820E-32
		x"0000000000000000000000000000000043429448190325000512000000000001291081", -- LUT(33) = log (1.000000000000000000000000000000010) = 4.3429448190325182765112891891660291082198748954452831046985920015492966E-33
		x"0000000000000000000000000000000004342944819032500051200000000000148650", -- LUT(34) = log (1.0000000000000000000000000000000010) = 4.3429448190325182765112891891660486514715605417775274054999432486346827E-34
		x"0000000000000000000000000000000000434294481903250005120000000000015069", -- LUT(35) = log (1.00000000000000000000000000000000010) = 4.3429448190325182765112891891660506057967291064107518355800783733561198E-35
		x"0000000000000000000000000000000000043429448190325000512000000000001506"); -- LUT(36) = log (1.000000000000000000000000000000000010) = 4.3429448190325182765112891891660506057967291064107518355800783733561198E-36

-- ====== FIN declaraci�n
-- declaracion de meomria de log para la parte de x<1

type mem_logSh_P is array (0 to 9) of STD_LOGIC_VECTOR (8*P+7 downto 0); 
type mem_logSh_N is array (0 to 9) of STD_LOGIC_VECTOR (8*P+7 downto 0); 

signal vlog_ShP: mem_LogSh_P;
signal vlog_ShN: mem_LogSh_N;
signal log_lut: std_logic_vector(8*P+7 downto 0); 
signal log_lut_sh: std_logic_vector(4*P+7 downto 0);

signal log_lut_optP, log_lut_optN, log_lut_opt: std_logic_vector(8*P+7 downto 0); 
signal log_lut_opt_sh: std_logic_vector(4*P+7 downto 0);

signal index:std_logic_vector(log2sup(2*P+1)-1 downto 0);

begin

	index <= (others => '0') when (conv_integer(true_step)>(P+2)) else true_step;


	vlog_ShP(0) <= (others => '0');
	vlog_ShP(1) <= lut_LogShP1(conv_integer(index));
	vlog_ShP(2) <= lut_LogShP2(conv_integer(index));
	vlog_ShP(3) <= lut_LogShP3(conv_integer(index));
	vlog_ShP(4) <= lut_LogShP4(conv_integer(index));
	vlog_ShP(5) <= lut_LogShP5(conv_integer(index));
	vlog_ShP(6) <= lut_LogShP6(conv_integer(index));
	vlog_ShP(7) <= lut_LogShP7(conv_integer(index));
	vlog_ShP(8) <= lut_LogShP8(conv_integer(index));
	vlog_ShP(9) <= lut_LogShP9(conv_integer(index));

	vlog_ShN(0) <= lut_LogShN0(conv_integer(index));
	vlog_ShN(1) <= lut_LogShN1(conv_integer(index));
	vlog_ShN(2) <= lut_LogShN2(conv_integer(index));
	vlog_ShN(3) <= lut_LogShN3(conv_integer(index));
	vlog_ShN(4) <= lut_LogShN4(conv_integer(index));
	vlog_ShN(5) <= lut_LogShN5(conv_integer(index));
	vlog_ShN(6) <= lut_LogShN6(conv_integer(index));
	vlog_ShN(7) <= lut_LogShN7(conv_integer(index));
	vlog_ShN(8) <= lut_LogShN8(conv_integer(index));
	vlog_ShN(9) <= lut_LogShN9(conv_integer(index));

	
	log_lut <= vlog_ShP(conv_integer(d)) when (x_greater_1='1') else vlog_ShN(conv_integer(d));

	
	log_lut_sh  <= log_lut(8*P+7 downto 4*P) when (offset_step="000000") else
					log_lut(8*P+3 downto 4*(P-1)) when (offset_step="000001") else
					log_lut(8*P-1 downto 4*(P-2)) when (offset_step="000010") else
					log_lut(8*P-5 downto 4*(P-3)) when (offset_step="000011") else
					log_lut(8*(P-1)-1 downto 4*(P-4)) when (offset_step="000100") else
					log_lut(8*(P-1)-5 downto 4*(P-5)) when (offset_step="000101") else
					log_lut(8*(P-2)-1 downto 4*(P-6)) when (offset_step="000110") else
					log_lut(8*(P-2)-5 downto 4*(P-7)) when (offset_step="000111") else
					log_lut(8*(P-3)-1 downto 4*(P-8)) when (offset_step="001000") else
					log_lut(8*(P-3)-5 downto 4*(P-9)) when (offset_step="001001") else
					log_lut(8*(P-4)-1 downto 4*(P-10)) when (offset_step="001010") else
					log_lut(8*(P-4)-5 downto 4*(P-11)) when (offset_step="001011") else
					log_lut(8*(P-5)-1 downto 4*(P-12)) when (offset_step="001100") else
					log_lut(8*(P-5)-5 downto 4*(P-13)) when (offset_step="001101") else
					log_lut(8*(P-6)-1 downto 4*(P-14)) when (offset_step="001110") else
					log_lut(8*(P-6)-5 downto 4*(P-15)) when (offset_step="001111") else
					log_lut(8*(P-7)-1 downto 4*(P-16)) when (offset_step="010000") else
					log_lut(8*(P-7)-5 downto 4*(P-17)) when (offset_step="010001") else
					log_lut(8*(P-8)-1 downto 4*(P-18)) when (offset_step="010010") else
					log_lut(8*(P-8)-5 downto 4*(P-19)) when (offset_step="010011") else
					log_lut(8*(P-9)-1 downto 4*(P-20)) when (offset_step="010100") else
					log_lut(8*(P-9)-5 downto 4*(P-21)) when (offset_step="010101") else
					log_lut(8*(P-10)-1 downto 4*(P-22)) when (offset_step="010110") else
					log_lut(8*(P-10)-5 downto 4*(P-23)) when (offset_step="010111") else
					log_lut(8*(P-11)-1 downto 4*(P-24)) when (offset_step="011000") else
					log_lut(8*(P-11)-5 downto 4*(P-25)) when (offset_step="011001") else
					log_lut(8*(P-12)-1 downto 4*(P-26)) when (offset_step="011010") else
					log_lut(8*(P-12)-5 downto 4*(P-27)) when (offset_step="011011") else
					log_lut(8*(P-13)-1 downto 4*(P-28)) when (offset_step="011100") else
					log_lut(8*(P-13)-5 downto 4*(P-29)) when (offset_step="011101") else
					log_lut(8*(P-14)-1 downto 4*(P-30)) when (offset_step="011110") else
					log_lut(8*(P-14)-5 downto 4*(P-31)) when (offset_step="011111") else
					log_lut(8*(P-15)-1 downto 4*(P-32)) when (offset_step="100000") else
					log_lut(8*(P-15)-5 downto 4*(P-33)) when (offset_step="100001") else
					log_lut(8*(P-16)-1 downto 4*(P-34)) when (offset_step="100010") else
					(others => '0');
	

	-- para LUT(P+2), se usa cuando hay 9's iniciales. 
	-- Lo que se debe hacer es desplazar a la derecha true_step - (P+2), por tema de patr�n
	-- y luego desplazar a la izquierda offset_step por tema de 9's iniciales. 
	-- Entonces desplazo a izquierda offset_step - true_step + P + 2. eso es igual a 
	-- P+2-step. Es decir que desplaza a P+2-step lugares a la izquierda Lut(P+2)
	
	log_lut_optP <= lut_LogShP1(P+2) when d=x"1" else
							lut_LogShP2(P+2) when d=x"2" else
							lut_LogShP3(P+2) when d=x"3" else
							lut_LogShP4(P+2) when d=x"4" else
							lut_LogShP5(P+2) when d=x"5" else
							lut_LogShP6(P+2) when d=x"6" else
							lut_LogShP7(P+2) when d=x"7" else
							lut_LogShP8(P+2) when d=x"8" else
							lut_LogShP9(P+2) when d=x"9" else
							(others => '0');
	
	log_lut_optN <= lut_LogShN0(P+2) when d=x"1" else
							lut_LogShN1(P+2) when d=x"1" else
							lut_LogShN2(P+2) when d=x"2" else
							lut_LogShN3(P+2) when d=x"3" else
							lut_LogShN4(P+2) when d=x"4" else
							lut_LogShN5(P+2) when d=x"5" else
							lut_LogShN6(P+2) when d=x"6" else
							lut_LogShN7(P+2) when d=x"7" else
							lut_LogShN8(P+2) when d=x"8" else
							lut_LogShN9(P+2) when d=x"9" else
							(others => '0');

	
	log_lut_opt <= log_lut_optP when (x_greater_1='1') else log_lut_optN;


	log_lut_opt_sh  <= log_lut_opt(4*(P+35)-1 downto 132) when (step="100011") else -- desplazo P-33 lugares a la izquierda  
							log_lut_opt(4*(P+34)-1 downto 128) when (step="100010") else -- desplazo P-32 lugares a la izquierda
							log_lut_opt(4*(P+33)-1 downto 124) when (step="100001") else -- desplazo P-31 lugares a la izquierda
							log_lut_opt(4*(P+32)-1 downto 120) when (step="100000") else -- desplazo P-30 lugares a la izquierda
							log_lut_opt(4*(P+31)-1 downto 116) when (step="011111") else
							log_lut_opt(4*(P+30)-1 downto 112) when (step="011110") else
							log_lut_opt(4*(P+29)-1 downto 108) when (step="011101") else
							log_lut_opt(4*(P+28)-1 downto 104) when (step="011100") else
							log_lut_opt(4*(P+27)-1 downto 100) when (step="011011") else
							log_lut_opt(4*(P+26)-1 downto 96) when (step="011010") else
							log_lut_opt(4*(P+25)-1 downto 92) when (step="011001") else
							log_lut_opt(4*(P+24)-1 downto 88) when (step="011000") else
							log_lut_opt(4*(P+23)-1 downto 84) when (step="010111") else
							log_lut_opt(4*(P+22)-1 downto 80) when (step="010110") else
							log_lut_opt(4*(P+21)-1 downto 76) when (step="010101") else
							log_lut_opt(4*(P+20)-1 downto 72) when (step="010100") else
							log_lut_opt(4*(P+19)-1 downto 68) when (step="010011") else
							log_lut_opt(4*(P+18)-1 downto 64) when (step="010010") else
							log_lut_opt(4*(P+17)-1 downto 60) when (step="010001") else
							log_lut_opt(4*(P+16)-1 downto 56) when (step="010000") else
							log_lut_opt(4*(P+15)-1 downto 52) when (step="001111") else
							log_lut_opt(4*(P+14)-1 downto 48) when (step="001110") else
							log_lut_opt(4*(P+13)-1 downto 44) when (step="001101") else
							log_lut_opt(4*(P+12)-1 downto 40) when (step="001100") else
							log_lut_opt(4*(P+11)-1 downto 36) when (step="001011") else
							log_lut_opt(4*(P+10)-1 downto 32) when (step="001010") else
							log_lut_opt(4*(P+9)-1 downto 28) when (step="001001") else
							log_lut_opt(4*(P+8)-1 downto 24) when (step="001000") else
							log_lut_opt(4*(P+7)-1 downto 20) when (step="000111") else
							log_lut_opt(4*(P+6)-1 downto 16) when (step="000110") else
							log_lut_opt(4*(P+5)-1 downto 12) when (step="000101") else
							log_lut_opt(4*(P+4)-1 downto 8) when (step="000100") else
							log_lut_opt(4*(P+3)-1 downto 4) when (step="000011") else
							log_lut_opt(4*(P+2)-1 downto 0) when (step="000010") else -- desplazo P lugares a la izquierda
							((log_lut_opt(4*(P+1)-1 downto 0))&(x"0")) when (step="000001") else -- desplazo P+1 lugares a la izquierda
							(others => '0');
	


	log(4*P+7 downto 0) <= log_lut_opt_sh when (conv_integer(true_step)>(P+2)) else log_lut_sh;
	log(4*P+8) <= x_greater_1;


end Behavioral;
